magic
tech sky130l
timestamp 1726446686
<< ndiffusion >>
rect 11 30 40 45
rect 11 22 18 30
rect 28 22 40 30
rect 11 16 40 22
rect 52 42 80 45
rect 52 28 63 42
rect 77 28 80 42
rect 52 16 80 28
<< ndc >>
rect 18 22 28 30
rect 63 28 77 42
<< ntransistor >>
rect 40 16 52 45
<< pdiffusion >>
rect 11 88 40 90
rect 11 80 18 88
rect 28 80 40 88
rect 11 61 40 80
rect 52 78 80 90
rect 52 64 63 78
rect 77 64 80 78
rect 52 61 80 64
<< pdc >>
rect 18 80 28 88
rect 63 64 77 78
<< ptransistor >>
rect 40 61 52 90
<< polysilicon >>
rect 40 90 52 95
rect 40 59 52 61
rect 1 47 52 59
rect 40 45 52 47
rect 40 11 52 16
<< m1 >>
rect 15 88 31 113
rect 15 80 18 88
rect 28 80 31 88
rect 15 77 31 80
rect 60 78 80 81
rect 60 64 63 78
rect 77 64 80 78
rect 60 59 80 64
rect 60 47 107 59
rect 60 42 80 47
rect 15 30 31 33
rect 15 22 18 30
rect 28 22 31 30
rect 60 28 63 42
rect 77 28 80 42
rect 60 26 80 28
rect 15 -3 31 22
<< labels >>
rlabel polysilicon 1 47 52 59 7 in
rlabel m1 60 47 107 59 3 out
rlabel m1 15 -3 31 22 5 GND!
rlabel m1 15 88 31 113 1 Vdd!
<< end >>
