magic
tech sky130l
timestamp 1734209687
<< ndiffusion >>
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 6 13 8
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 8 12 11
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 28 13 29
rect 8 25 9 28
rect 12 25 13 28
rect 8 19 13 25
rect 15 24 20 29
rect 15 21 16 24
rect 19 21 20 24
rect 15 19 20 21
<< pdc >>
rect 9 25 12 28
rect 16 21 19 24
<< ptransistor >>
rect 13 19 15 29
<< polysilicon >>
rect 13 29 15 31
rect 13 17 15 19
rect 23 18 28 19
rect 23 17 24 18
rect 13 15 24 17
rect 27 15 28 18
rect 13 12 15 15
rect 23 14 28 15
rect 13 4 15 6
<< pc >>
rect 24 15 27 18
<< m1 >>
rect 8 35 12 36
rect 8 32 9 35
rect 9 28 12 32
rect 9 24 12 25
rect 15 21 16 24
rect 19 21 23 24
rect 26 21 27 24
rect 16 15 24 18
rect 27 15 28 18
rect 9 11 12 12
rect 8 8 9 9
rect 16 11 19 15
rect 12 8 13 9
rect 8 7 13 8
rect 16 7 19 8
rect 6 4 13 7
rect 6 3 12 4
rect 24 0 28 8
<< m2c >>
rect 9 32 12 35
rect 23 21 26 24
rect 9 8 12 11
rect 24 8 27 11
<< m2 >>
rect 8 35 13 36
rect 8 32 9 35
rect 12 32 13 35
rect 8 31 13 32
rect 22 24 27 25
rect 22 21 23 24
rect 26 21 27 24
rect 22 20 27 21
rect 23 12 25 20
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 7 13 8
rect 23 11 28 12
rect 23 8 24 11
rect 27 8 28 11
rect 23 7 28 8
rect 6 4 13 7
rect 6 3 12 4
<< labels >>
rlabel pdiffusion 16 20 16 20 3 Y
rlabel polysilicon 14 13 14 13 3 x
rlabel polysilicon 14 18 14 18 3 x
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 25 5 25 5 3 Y
port 2 e
rlabel m2 8 35 13 36 4 Vdd
rlabel m2 8 4 13 8 2 GND
<< end >>
