magic
tech sky130l
timestamp 1731041890
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
<< pdiffusion >>
rect 8 23 13 34
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 19 20 34
rect 22 33 27 34
rect 22 30 23 33
rect 26 30 27 33
rect 22 19 27 30
<< pdc >>
rect 9 20 12 23
rect 23 30 26 33
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
<< polysilicon >>
rect 15 44 20 45
rect 15 42 16 44
rect 13 41 16 42
rect 19 41 20 44
rect 13 40 20 41
rect 13 34 15 40
rect 20 34 22 36
rect 30 34 35 35
rect 30 31 31 34
rect 34 31 35 34
rect 30 30 35 31
rect 13 12 15 19
rect 20 17 22 19
rect 32 17 34 30
rect 20 15 34 17
rect 20 12 22 15
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 16 41 19 44
rect 31 31 34 34
<< m1 >>
rect 16 44 20 45
rect 19 41 20 44
rect 16 36 20 41
rect 24 44 28 45
rect 27 41 28 44
rect 24 39 28 41
rect 32 39 36 45
rect 23 36 28 39
rect 31 36 36 39
rect 23 33 26 36
rect 31 34 34 36
rect 31 30 34 31
rect 23 29 26 30
rect 9 23 12 24
rect 9 16 12 20
rect 9 13 26 16
rect 9 10 12 13
rect 23 10 26 13
rect 8 7 9 8
rect 15 7 16 10
rect 19 7 20 10
rect 8 4 12 7
rect 23 6 26 7
rect 35 5 36 8
rect 32 4 36 5
<< m2c >>
rect 24 41 27 44
rect 16 7 19 10
rect 32 5 35 8
<< m2 >>
rect 23 44 28 45
rect 23 41 24 44
rect 27 41 28 44
rect 23 40 28 41
rect 15 10 20 11
rect 15 7 16 10
rect 19 9 34 10
rect 19 8 36 9
rect 19 7 20 8
rect 15 6 20 7
rect 31 5 32 8
rect 35 5 36 8
rect 31 4 36 5
<< labels >>
rlabel polysilicon 21 13 21 13 3 B
rlabel polysilicon 21 18 21 18 3 B
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel m1 9 5 9 5 3 Y
port 4 e
rlabel m1 33 37 33 37 3 B
port 3 e
rlabel m1 17 37 17 37 3 A
port 5 e
rlabel m1 33 5 33 5 3 GND
port 1 e
rlabel m2 27 40 28 45 5 Vdd
<< end >>
