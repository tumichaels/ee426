magic
tech sky130l
timestamp 1726535576
<< rotate >>
rect 94 185 142 190
<< polysilicon >>
rect 13 77 32 82
rect 103 77 122 82
rect 13 61 32 66
rect 103 61 122 66
rect 13 24 32 29
rect 103 24 122 29
rect 13 8 32 13
rect 103 8 122 13
<< pc >>
rect 46 262 54 268
rect 79 186 82 189
rect 95 186 98 189
<< m1 >>
rect 44 320 56 366
rect -4 201 9 284
rect 44 268 56 270
rect 44 262 46 268
rect 54 262 56 268
rect 44 224 56 262
rect 92 245 103 284
rect 156 245 166 246
rect 92 241 166 245
rect 101 238 166 241
rect 44 217 76 224
rect -4 196 105 201
rect -4 158 9 196
rect 45 189 83 190
rect 45 186 79 189
rect 82 186 83 189
rect 45 185 83 186
rect 94 189 142 190
rect 94 186 95 189
rect 98 186 142 189
rect 94 185 142 186
rect 24 158 31 159
rect -4 153 31 158
rect 24 142 31 153
rect 45 146 52 185
rect 135 145 142 185
rect 156 112 166 238
rect 8 -10 20 -8
rect 8 -14 11 -10
rect 16 -14 20 -10
rect 8 -16 20 -14
rect 24 -37 31 42
rect 66 -10 73 2
rect 66 -13 68 -10
rect 71 -13 73 -10
rect 66 -15 73 -13
rect 114 -37 121 41
rect 156 -10 163 3
rect 156 -13 158 -10
rect 161 -13 163 -10
rect 156 -14 163 -13
rect 10 -46 122 -37
rect 114 -47 121 -46
<< m2c >>
rect 11 -14 16 -10
rect 68 -13 71 -10
rect 158 -13 161 -10
<< m2 >>
rect 9 -10 163 -8
rect 9 -14 11 -10
rect 16 -13 68 -10
rect 71 -13 158 -10
rect 161 -13 163 -10
rect 16 -14 163 -13
rect 9 -16 163 -14
use inv  inv_0
timestamp 1726446686
transform 0 -1 103 1 0 259
box 1 -3 107 113
use nor2  nor2_0 ../nor
timestamp 1726527990
transform 0 -1 261 1 0 -71
box 256 151 316 194
use or4  or4_1
timestamp 1726533950
transform 1 0 148 0 1 -27
box -45 24 15 174
use or4  or4_0
timestamp 1726533950
transform 1 0 58 0 1 -27
box -45 24 15 174
<< labels >>
rlabel m2 9 -16 11 -8 7 GND!
rlabel m1 10 -46 122 -37 7 Vdd!
rlabel m1 44 320 56 366 1 out
rlabel polysilicon 13 77 32 82 7 in000
rlabel polysilicon 13 61 32 66 7 in001
rlabel polysilicon 13 24 32 29 7 in010
rlabel polysilicon 13 8 32 13 7 in011
rlabel polysilicon 103 77 122 82 7 in100
rlabel polysilicon 103 61 122 66 7 in101
rlabel polysilicon 103 24 122 29 7 in110
rlabel polysilicon 103 8 122 13 7 in111
<< end >>
