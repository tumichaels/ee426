magic
tech sky130l
timestamp 1734213373
<< ndiffusion >>
rect 8 15 13 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 10 13 12
rect 15 15 20 16
rect 15 12 16 15
rect 19 12 20 15
rect 15 10 20 12
rect 22 14 27 16
rect 22 11 23 14
rect 26 11 27 14
rect 22 10 27 11
rect 33 10 38 16
rect 33 7 34 10
rect 37 7 38 10
rect 33 6 38 7
rect 40 15 45 16
rect 40 12 41 15
rect 44 12 45 15
rect 40 6 45 12
rect 47 15 52 16
rect 47 12 48 15
rect 51 12 52 15
rect 47 6 52 12
rect 58 10 63 16
rect 58 7 59 10
rect 62 7 63 10
rect 58 6 63 7
rect 65 10 70 16
rect 65 7 66 10
rect 69 7 70 10
rect 65 6 70 7
rect 72 15 77 16
rect 72 12 73 15
rect 76 12 77 15
rect 72 6 77 12
<< ndc >>
rect 9 12 12 15
rect 16 12 19 15
rect 23 11 26 14
rect 34 7 37 10
rect 41 12 44 15
rect 48 12 51 15
rect 59 7 62 10
rect 66 7 69 10
rect 73 12 76 15
<< ntransistor >>
rect 13 10 15 16
rect 20 10 22 16
rect 38 6 40 16
rect 45 6 47 16
rect 63 6 65 16
rect 70 6 72 16
<< pdiffusion >>
rect 8 27 13 31
rect 8 24 9 27
rect 12 24 13 27
rect 8 23 13 24
rect 15 30 20 31
rect 15 27 16 30
rect 19 27 20 30
rect 15 23 20 27
rect 22 27 27 31
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 33 27 38 38
rect 33 24 34 27
rect 37 24 38 27
rect 33 23 38 24
rect 40 27 45 38
rect 40 24 41 27
rect 44 24 45 27
rect 40 23 45 24
rect 47 27 52 38
rect 47 24 48 27
rect 51 24 52 27
rect 47 23 52 24
rect 58 27 63 38
rect 58 24 59 27
rect 62 24 63 27
rect 58 23 63 24
rect 65 37 70 38
rect 65 34 66 37
rect 69 34 70 37
rect 65 23 70 34
rect 72 27 77 38
rect 72 24 73 27
rect 76 24 77 27
rect 72 23 77 24
<< pdc >>
rect 9 24 12 27
rect 16 27 19 30
rect 23 24 26 27
rect 34 24 37 27
rect 41 24 44 27
rect 48 24 51 27
rect 59 24 62 27
rect 66 34 69 37
rect 73 24 76 27
<< ptransistor >>
rect 13 23 15 31
rect 20 23 22 31
rect 38 23 40 38
rect 45 23 47 38
rect 63 23 65 38
rect 70 23 72 38
<< polysilicon >>
rect 62 45 67 46
rect 25 43 30 44
rect 25 40 26 43
rect 29 42 30 43
rect 62 42 63 45
rect 66 42 67 45
rect 75 45 80 46
rect 75 42 76 45
rect 79 42 80 45
rect 29 40 40 42
rect 62 41 67 42
rect 70 41 80 42
rect 25 39 30 40
rect 10 38 15 39
rect 38 38 40 40
rect 45 38 47 40
rect 63 38 65 41
rect 70 40 77 41
rect 70 38 72 40
rect 10 35 11 38
rect 14 35 15 38
rect 10 34 15 35
rect 13 31 15 34
rect 20 31 22 33
rect 13 16 15 23
rect 20 20 22 23
rect 38 20 40 23
rect 20 18 40 20
rect 20 16 22 18
rect 38 16 40 18
rect 45 16 47 23
rect 63 16 65 23
rect 70 16 72 23
rect 13 8 15 10
rect 20 8 22 10
rect 25 6 30 7
rect 25 3 26 6
rect 29 3 30 6
rect 38 4 40 6
rect 25 2 30 3
rect 28 1 30 2
rect 45 1 47 6
rect 63 4 65 6
rect 70 4 72 6
rect 28 -1 47 1
<< pc >>
rect 26 40 29 43
rect 63 42 66 45
rect 76 42 79 45
rect 11 35 14 38
rect 26 3 29 6
<< m1 >>
rect 8 40 14 51
rect 29 44 35 51
rect 44 49 53 51
rect 44 46 48 49
rect 51 46 53 49
rect 44 45 53 46
rect 63 45 66 46
rect 76 45 79 46
rect 25 43 36 44
rect 25 40 26 43
rect 29 40 36 43
rect 11 38 14 40
rect 48 37 51 45
rect 66 42 67 45
rect 63 41 66 42
rect 56 37 59 38
rect 11 34 14 35
rect 17 34 66 37
rect 69 34 70 37
rect 76 36 79 42
rect 17 31 20 34
rect 16 30 20 31
rect 9 27 12 28
rect 19 28 20 30
rect 16 26 19 27
rect 23 27 26 28
rect 41 27 44 28
rect 9 15 12 24
rect 33 24 34 27
rect 37 24 38 27
rect 47 24 48 27
rect 51 24 59 27
rect 62 24 63 27
rect 72 24 73 27
rect 76 24 77 27
rect 9 11 12 12
rect 16 15 19 16
rect 16 11 19 12
rect 23 14 26 24
rect 41 15 44 24
rect 49 16 75 18
rect 48 15 75 16
rect 26 11 29 13
rect 40 12 41 15
rect 44 12 45 15
rect 51 12 52 15
rect 72 12 73 15
rect 76 12 77 15
rect 48 11 51 12
rect 23 10 29 11
rect 8 7 9 8
rect 6 6 9 7
rect 4 5 9 6
rect 4 2 12 5
rect 26 6 29 10
rect 34 10 37 11
rect 66 10 69 11
rect 37 8 40 9
rect 55 8 59 10
rect 37 7 59 8
rect 62 7 63 10
rect 69 7 77 9
rect 34 6 58 7
rect 66 6 77 7
rect 80 8 83 9
rect 80 6 84 8
rect 37 5 58 6
rect 26 2 29 3
rect 4 -2 11 2
rect 77 -1 84 6
<< m2c >>
rect 48 46 51 49
rect 11 35 14 38
rect 67 42 70 45
rect 76 33 79 36
rect 9 24 12 27
rect 34 24 37 27
rect 16 12 19 15
rect 41 12 44 15
rect 9 5 12 8
rect 77 6 80 9
<< m2 >>
rect 44 49 53 51
rect 44 46 48 49
rect 51 46 53 49
rect 44 45 53 46
rect 66 45 71 46
rect 66 42 67 45
rect 70 42 71 45
rect 66 41 71 42
rect 10 38 15 39
rect 10 35 11 38
rect 14 36 15 38
rect 67 36 69 41
rect 14 35 69 36
rect 10 34 69 35
rect 75 36 80 37
rect 75 33 76 36
rect 79 33 80 36
rect 75 32 80 33
rect 29 31 42 32
rect 64 31 78 32
rect 11 30 78 31
rect 11 29 31 30
rect 40 29 66 30
rect 11 28 13 29
rect 8 27 13 28
rect 8 24 9 27
rect 12 24 13 27
rect 8 23 13 24
rect 33 27 38 28
rect 72 27 77 28
rect 33 24 34 27
rect 37 25 77 27
rect 37 24 38 25
rect 33 23 38 24
rect 72 23 77 25
rect 36 18 69 20
rect 36 16 38 18
rect 15 15 38 16
rect 15 12 16 15
rect 19 14 38 15
rect 40 15 45 16
rect 19 12 20 14
rect 15 11 20 12
rect 40 12 41 15
rect 44 12 45 15
rect 40 11 45 12
rect 40 9 42 11
rect 8 8 42 9
rect 8 5 9 8
rect 12 7 42 8
rect 67 9 69 18
rect 76 9 81 10
rect 67 7 77 9
rect 12 5 13 7
rect 76 6 77 7
rect 80 8 81 9
rect 80 6 84 8
rect 76 5 84 6
rect 8 4 13 5
rect 77 -1 84 5
<< labels >>
rlabel m1 8 40 12 44 4 B
rlabel m1 32 40 36 44 5 A
rlabel m1 6 2 12 5 2 Y
rlabel m2 44 45 48 51 5 Vdd
rlabel m2 80 4 84 8 7 GND
<< end >>
