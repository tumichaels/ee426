magic
tech TSMC180
timestamp 1734149807
<< ndiffusion >>
rect 6 10 12 12
rect 6 8 7 10
rect 9 8 12 10
rect 6 7 12 8
rect 14 11 20 12
rect 14 9 16 11
rect 18 9 20 11
rect 14 7 20 9
rect 22 11 28 12
rect 22 9 24 11
rect 26 9 28 11
rect 22 7 28 9
rect 30 11 36 12
rect 30 9 33 11
rect 35 9 36 11
rect 30 7 36 9
<< ndcontact >>
rect 7 8 9 10
rect 16 9 18 11
rect 24 9 26 11
rect 33 9 35 11
<< ntransistor >>
rect 12 7 14 12
rect 20 7 22 12
rect 28 7 30 12
<< pdiffusion >>
rect 6 31 12 43
rect 6 29 8 31
rect 10 29 12 31
rect 6 28 12 29
rect 14 28 20 43
rect 22 42 26 43
rect 22 40 23 42
rect 25 40 26 42
rect 22 36 26 40
rect 22 28 28 36
rect 30 31 36 36
rect 30 29 33 31
rect 35 29 36 31
rect 30 28 36 29
<< pdcontact >>
rect 8 29 10 31
rect 23 40 25 42
rect 33 29 35 31
<< ptransistor >>
rect 12 28 14 43
rect 20 28 22 43
rect 28 28 30 36
<< polysilicon >>
rect 10 49 14 50
rect 10 47 11 49
rect 13 47 14 49
rect 10 46 14 47
rect 18 49 22 50
rect 18 47 19 49
rect 21 47 22 49
rect 18 46 22 47
rect 12 43 14 46
rect 20 43 22 46
rect 28 36 30 39
rect 12 12 14 28
rect 20 12 22 28
rect 28 23 30 28
rect 28 22 32 23
rect 28 20 29 22
rect 31 20 32 22
rect 28 19 32 20
rect 28 12 30 19
rect 12 4 14 7
rect 20 4 22 7
rect 28 4 30 7
<< polycontact >>
rect 11 47 13 49
rect 19 47 21 49
rect 29 20 31 22
<< m1 >>
rect 6 50 9 57
rect 22 50 25 57
rect 6 49 14 50
rect 6 47 11 49
rect 13 47 14 49
rect 10 46 14 47
rect 18 49 25 50
rect 18 47 19 49
rect 21 47 25 49
rect 18 46 22 47
rect 33 43 36 57
rect 22 42 36 43
rect 22 40 23 42
rect 25 40 36 42
rect 22 39 26 40
rect 7 31 11 32
rect 7 29 8 31
rect 10 29 11 31
rect 7 28 11 29
rect 32 31 40 32
rect 32 29 33 31
rect 35 29 40 31
rect 32 28 40 29
rect 8 22 11 28
rect 28 22 32 23
rect 8 20 29 22
rect 31 20 32 22
rect 8 19 32 20
rect 16 12 19 19
rect 37 12 40 28
rect 15 11 19 12
rect 6 10 10 11
rect 6 8 7 10
rect 9 8 10 10
rect 15 9 16 11
rect 18 9 19 11
rect 15 8 19 9
rect 23 11 27 12
rect 23 9 24 11
rect 26 9 27 11
rect 23 8 27 9
rect 32 11 40 12
rect 32 9 33 11
rect 35 9 40 11
rect 32 8 40 9
rect 6 5 10 8
rect 23 5 26 8
rect 6 2 26 5
rect 6 -3 9 2
rect 37 -3 40 8
<< labels >>
rlabel pdiffusion 31 29 31 29 3 Y
rlabel ndiffusion 31 8 31 8 3 Y
rlabel polysilicon 29 13 29 13 3 _Y
rlabel polysilicon 29 26 29 26 3 _Y
rlabel ndiffusion 23 8 23 8 3 GND
rlabel pdiffusion 23 29 23 29 3 Vdd
rlabel polysilicon 21 13 21 13 3 A
rlabel polysilicon 21 26 21 26 3 A
rlabel ndiffusion 15 8 15 8 3 _Y
rlabel polysilicon 13 13 13 13 3 B
rlabel polysilicon 13 26 13 26 3 B
rlabel ndiffusion 7 8 7 8 3 GND
rlabel pdiffusion 7 29 7 29 3 _Y
rlabel m1 19 48 19 48 3 A
port 5 e
rlabel m1 7 48 7 48 3 B
port 3 e
rlabel m1 7 11 7 11 3 GND
port 1 e
rlabel m1 38 30 38 30 3 Y
port 4 e
rlabel m1 34 48 34 48 3 Vdd
port 2 e
<< end >>
