magic
tech sky130l
timestamp 1726582099
<< polysilicon >>
rect 1 159 19 160
rect 1 156 3 159
rect 6 156 19 159
rect 1 155 19 156
rect -9 143 19 144
rect -9 140 -7 143
rect -4 140 19 143
rect -9 139 19 140
rect -19 91 19 96
rect -19 75 19 80
rect -19 27 19 32
rect -19 11 19 16
<< pc >>
rect 3 156 6 159
rect -7 140 -4 143
<< m1 >>
rect 1 159 8 160
rect 1 156 3 159
rect 6 156 8 159
rect -9 143 -2 144
rect -9 140 -7 143
rect -4 140 -2 143
rect -9 56 -2 140
rect 1 120 8 156
rect 1 115 2 120
rect 7 115 8 120
rect 1 114 8 115
rect -9 51 -8 56
rect -3 51 -2 56
rect -9 50 -2 51
rect 11 -10 18 171
rect 32 160 39 171
rect 32 120 39 121
rect 32 115 33 120
rect 38 115 39 120
rect 32 107 39 115
rect 32 56 39 57
rect 32 51 33 56
rect 38 51 39 56
rect 32 43 39 51
rect 53 -10 60 171
<< m2c >>
rect 2 115 7 120
rect -8 51 -3 56
rect 33 115 38 120
rect 33 51 38 56
<< m2 >>
rect 1 120 39 121
rect 1 115 2 120
rect 7 115 33 120
rect 38 115 39 120
rect 1 114 39 115
rect -9 56 39 57
rect -9 51 -8 56
rect -3 51 33 56
rect 38 51 39 56
rect -9 50 39 51
use nand2  nand2_0 ../nand
timestamp 1726527220
transform 1 0 -44 0 1 97
box 44 31 104 74
use nor2  nor2_1
timestamp 1726527990
transform 1 0 -256 0 1 -87
box 256 151 316 194
use nor2  nor2_0
timestamp 1726527990
transform 1 0 -256 0 1 -151
box 256 151 316 194
<< labels >>
rlabel m1 11 -10 18 171 5 Vdd!
rlabel m1 53 -10 60 171 5 GND!
rlabel m1 32 160 39 171 1 out
rlabel polysilicon -19 91 19 96 7 in00
rlabel polysilicon -19 75 19 80 7 in01
rlabel polysilicon -19 27 19 32 7 in10
rlabel polysilicon -19 11 19 16 7 in11
<< end >>
