magic
tech sky130l
timestamp 1729862358
<< ndiffusion >>
rect 8 15 13 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 10 13 12
rect 41 10 44 16
rect 46 15 53 16
rect 46 12 48 15
rect 51 12 53 15
rect 46 10 53 12
rect 49 8 53 10
rect 55 8 58 16
rect 60 15 65 16
rect 60 12 61 15
rect 64 12 65 15
rect 60 10 65 12
rect 69 15 74 16
rect 69 12 70 15
rect 73 12 74 15
rect 69 10 74 12
rect 60 8 64 10
<< ndc >>
rect 9 12 12 15
rect 48 12 51 15
rect 61 12 64 15
rect 70 12 73 15
<< ntransistor >>
rect 13 10 41 16
rect 44 10 46 16
rect 53 8 55 16
rect 58 8 60 16
rect 65 10 69 16
<< pdiffusion >>
rect 49 29 53 34
rect 8 27 13 29
rect 8 24 9 27
rect 12 24 13 27
rect 8 23 13 24
rect 27 23 44 29
rect 46 27 53 29
rect 46 24 48 27
rect 51 24 53 27
rect 46 23 53 24
rect 55 23 58 34
rect 60 33 64 34
rect 60 27 65 33
rect 60 24 61 27
rect 64 24 65 27
rect 60 23 65 24
rect 69 27 74 33
rect 69 24 70 27
rect 73 24 74 27
rect 69 23 74 24
<< pdc >>
rect 9 24 12 27
rect 48 24 51 27
rect 61 24 64 27
rect 70 24 73 27
<< ptransistor >>
rect 13 23 27 29
rect 44 23 46 29
rect 53 23 55 34
rect 58 23 60 34
rect 65 23 69 33
<< polysilicon >>
rect 36 39 55 40
rect 24 38 29 39
rect 16 36 21 37
rect 16 33 17 36
rect 20 33 21 36
rect 24 35 25 38
rect 28 36 29 38
rect 36 36 37 39
rect 40 38 55 39
rect 40 36 41 38
rect 51 36 55 38
rect 28 35 32 36
rect 36 35 41 36
rect 24 34 32 35
rect 53 34 55 36
rect 58 34 60 37
rect 16 31 21 33
rect 30 32 32 34
rect 13 29 27 31
rect 30 30 46 32
rect 44 29 46 30
rect 65 33 69 35
rect 13 21 27 23
rect 13 16 41 18
rect 44 16 46 23
rect 53 16 55 23
rect 58 16 60 23
rect 65 21 69 23
rect 77 21 82 22
rect 65 18 78 21
rect 81 18 82 21
rect 65 16 69 18
rect 77 17 82 18
rect 13 8 41 10
rect 44 8 46 10
rect 65 8 69 10
rect 53 4 55 8
rect 58 4 60 8
<< pc >>
rect 17 33 20 36
rect 25 35 28 38
rect 37 36 40 39
rect 78 18 81 21
<< m1 >>
rect 8 36 12 40
rect 32 39 36 40
rect 24 38 29 39
rect 16 36 21 37
rect 16 33 17 36
rect 20 33 21 36
rect 24 35 25 38
rect 28 35 29 38
rect 32 36 37 39
rect 40 36 41 39
rect 56 36 60 40
rect 80 36 84 40
rect 24 34 29 35
rect 16 32 21 33
rect 26 33 29 34
rect 79 35 84 36
rect 26 30 73 33
rect 79 32 80 35
rect 83 32 84 35
rect 69 28 73 30
rect 69 27 74 28
rect 8 24 9 27
rect 12 24 13 27
rect 47 24 48 27
rect 51 24 52 27
rect 60 24 61 27
rect 64 24 65 27
rect 69 24 70 27
rect 73 24 74 27
rect 8 15 13 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 11 13 12
rect 48 15 51 24
rect 69 23 74 24
rect 70 16 73 23
rect 78 21 81 22
rect 60 15 65 16
rect 60 12 61 15
rect 64 12 65 15
rect 69 15 74 16
rect 69 12 70 15
rect 73 12 74 15
rect 48 8 51 12
rect 78 8 81 18
rect 8 5 81 8
rect 8 4 12 5
<< m2c >>
rect 80 32 83 35
rect 9 24 12 27
rect 61 24 64 27
rect 9 12 12 15
rect 61 12 64 15
<< m2 >>
rect 79 35 84 36
rect 79 32 80 35
rect 83 32 84 35
rect 79 31 84 32
rect 8 27 13 28
rect 60 27 65 28
rect 8 24 9 27
rect 12 24 61 27
rect 64 24 65 27
rect 8 23 13 24
rect 60 23 65 24
rect 8 15 13 16
rect 60 15 65 16
rect 80 15 83 31
rect 8 12 9 15
rect 12 12 61 15
rect 64 12 83 15
rect 8 11 13 12
rect 60 11 65 12
<< m3pin >>
rect 9 12 12 15
<< labels >>
rlabel pdiffusion 70 24 70 24 3 #7
rlabel polysilicon 66 17 66 17 3 out
rlabel polysilicon 66 22 66 22 3 out
rlabel ndiffusion 70 11 70 11 3 #7
rlabel pdiffusion 61 24 61 24 3 Vdd
rlabel polysilicon 59 17 59 17 3 in(0)
rlabel polysilicon 59 22 59 22 3 in(0)
rlabel polysilicon 54 17 54 17 3 in(1)
rlabel polysilicon 54 22 54 22 3 in(1)
rlabel pdiffusion 47 24 47 24 3 out
rlabel polysilicon 45 17 45 17 3 #7
rlabel polysilicon 45 22 45 22 3 #7
rlabel polysilicon 14 17 14 17 3 Vdd
rlabel polysilicon 14 22 14 22 3 GND
rlabel ndiffusion 9 11 9 11 3 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m1 81 37 81 37 3 GND
port 1 e
rlabel m1 57 37 57 37 3 Vdd
port 2 e
rlabel m1 33 37 33 37 3 in(1)
port 3 e
rlabel m1 9 5 9 5 3 out
port 4 e
rlabel m1 9 37 9 37 3 in(0)
port 5 e
rlabel m1 50 11 50 11 1 out
rlabel m2 61 13 61 13 1 GND
<< end >>
