magic
tech sky130l
timestamp 1731020590
<< ndiffusion >>
rect 8 15 14 16
rect 8 12 9 15
rect 12 12 14 15
rect 8 6 14 12
rect 16 6 21 16
rect 23 14 28 16
rect 23 11 24 14
rect 27 11 28 14
rect 23 10 28 11
rect 30 15 36 16
rect 30 12 31 15
rect 35 12 36 15
rect 30 10 36 12
rect 23 6 27 10
<< ndc >>
rect 9 12 12 15
rect 24 11 27 14
rect 31 12 35 15
<< ntransistor >>
rect 14 6 16 16
rect 21 6 23 16
rect 28 10 30 16
<< pdiffusion >>
rect 8 30 14 31
rect 8 27 9 30
rect 12 27 14 30
rect 8 23 14 27
rect 16 28 21 31
rect 16 25 17 28
rect 20 25 21 28
rect 16 23 21 25
rect 23 30 28 31
rect 23 27 24 30
rect 27 27 28 30
rect 23 23 28 27
rect 30 30 36 31
rect 30 27 31 30
rect 35 27 36 30
rect 30 23 36 27
<< pdc >>
rect 9 27 12 30
rect 17 25 20 28
rect 24 27 27 30
rect 31 27 35 30
<< ptransistor >>
rect 14 23 16 31
rect 21 23 23 31
rect 28 23 30 31
<< polysilicon >>
rect 8 43 16 44
rect 8 40 9 43
rect 12 40 16 43
rect 8 39 16 40
rect 14 31 16 39
rect 21 43 28 44
rect 21 40 24 43
rect 27 40 28 43
rect 21 39 28 40
rect 21 31 23 39
rect 28 31 30 35
rect 14 16 16 23
rect 21 16 23 23
rect 28 16 30 23
rect 14 4 16 6
rect 21 4 23 6
rect 28 5 30 10
rect 28 4 36 5
rect 28 1 32 4
rect 35 1 36 4
rect 28 0 36 1
<< pc >>
rect 9 40 12 43
rect 24 40 27 43
rect 32 1 35 4
<< m1 >>
rect 19 45 20 48
rect 4 43 13 44
rect 4 40 9 43
rect 12 40 13 43
rect 4 39 13 40
rect 16 35 20 45
rect 24 44 28 48
rect 23 43 28 44
rect 23 40 24 43
rect 27 40 28 43
rect 23 39 28 40
rect 8 32 28 35
rect 8 30 13 32
rect 8 27 9 30
rect 12 27 13 30
rect 23 30 28 32
rect 32 31 36 48
rect 8 26 13 27
rect 16 28 20 29
rect 16 25 17 28
rect 23 27 24 30
rect 27 27 28 30
rect 23 26 28 27
rect 31 30 36 31
rect 35 27 36 30
rect 16 23 20 25
rect 16 22 24 23
rect 8 19 20 22
rect 23 19 24 22
rect 8 18 24 19
rect 8 15 13 18
rect 31 16 36 27
rect 30 15 36 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 11 13 12
rect 23 14 27 15
rect 23 11 24 14
rect 30 12 31 15
rect 35 12 36 15
rect 23 10 27 11
rect 8 1 9 4
rect 24 3 27 10
rect 12 1 27 3
rect 8 0 27 1
rect 31 8 36 9
rect 31 5 32 8
rect 35 5 36 8
rect 31 4 36 5
rect 31 1 32 4
rect 35 1 36 4
rect 31 0 36 1
<< m2c >>
rect 16 45 19 48
rect 20 19 23 22
rect 9 1 12 4
rect 32 5 35 8
<< m2 >>
rect 15 48 20 49
rect 15 45 16 48
rect 19 45 20 48
rect 15 44 20 45
rect 19 22 36 23
rect 19 19 20 22
rect 23 19 36 22
rect 19 18 36 19
rect 31 8 36 18
rect 31 5 32 8
rect 35 5 36 8
rect 8 4 13 5
rect 31 4 36 5
rect 8 1 9 4
rect 12 1 13 4
rect 8 0 13 1
<< labels >>
rlabel polysilicon 29 17 29 17 3 _Y
rlabel ndiffusion 31 11 31 11 3 Y
rlabel ndiffusion 10 7 10 7 3 _Y
rlabel pdiffusion 10 24 10 24 3 Vdd
rlabel pdiffusion 17 24 17 24 3 _Y
rlabel pdiffusion 24 24 24 24 3 Vdd
rlabel polysilicon 29 22 29 22 3 _Y
rlabel pdiffusion 31 24 31 24 3 Y
rlabel m1 17 45 17 45 3 Vdd
port 3 e
rlabel ndiffusion 24 7 24 7 3 GND
rlabel m1 9 1 9 1 3 GND
port 4 e
rlabel m1 33 45 33 45 3 Y
port 1 e
rlabel m1 4 39 9 44 3 A
rlabel m1 25 45 25 45 3 B
port 2 e
<< end >>
