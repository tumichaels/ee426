magic
tech sky130l
timestamp 1731046771
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
<< pdiffusion >>
rect 8 23 13 34
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 19 20 34
rect 22 33 27 34
rect 22 30 23 33
rect 26 30 27 33
rect 22 19 27 30
<< pdc >>
rect 9 20 12 23
rect 23 30 26 33
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
<< polysilicon >>
rect 9 45 15 46
rect 9 42 10 45
rect 13 42 15 45
rect 33 44 38 45
rect 33 42 34 44
rect 9 41 15 42
rect 13 34 15 41
rect 32 41 34 42
rect 37 41 38 44
rect 32 40 38 41
rect 20 34 22 36
rect 13 12 15 19
rect 20 17 22 19
rect 32 17 34 40
rect 20 15 34 17
rect 20 12 22 15
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 10 42 13 45
rect 34 41 37 44
<< m1 >>
rect 8 47 12 48
rect 8 45 13 47
rect 8 44 10 45
rect 10 41 13 42
rect 23 44 26 48
rect 32 44 39 48
rect 32 42 34 44
rect 23 33 26 41
rect 37 42 39 44
rect 34 40 37 41
rect 23 29 26 30
rect 9 23 12 24
rect 9 16 12 20
rect 9 13 26 16
rect 9 10 12 13
rect 23 10 26 13
rect 6 7 9 8
rect 15 7 16 10
rect 19 7 20 10
rect 6 2 12 7
rect 23 6 26 7
rect 35 5 36 8
rect 32 4 36 5
<< m2c >>
rect 23 41 26 44
rect 16 7 19 10
rect 32 5 35 8
<< m2 >>
rect 22 44 27 48
rect 22 41 23 44
rect 26 41 27 44
rect 22 40 27 41
rect 18 14 33 17
rect 18 11 20 14
rect 15 10 20 11
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
rect 31 9 33 14
rect 31 8 36 9
rect 31 5 32 8
rect 35 5 36 8
rect 31 4 36 5
<< labels >>
rlabel polysilicon 21 13 21 13 3 B
rlabel polysilicon 21 18 21 18 3 B
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel m1 9 5 9 5 3 Y
port 4 e
rlabel m1 33 5 33 5 3 GND
port 1 e
rlabel m1 8 44 12 48 5 A
rlabel m2 22 44 27 48 5 Vdd
rlabel m1 32 42 39 48 6 B
<< end >>
