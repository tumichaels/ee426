magic
tech sky130l
timestamp 0
<< end >>
