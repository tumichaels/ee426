magic
tech sky130l
timestamp 1731040958
<< ndiffusion >>
rect 8 15 13 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 10 13 12
rect 41 10 44 16
rect 46 15 53 16
rect 46 12 48 15
rect 51 12 53 15
rect 46 10 53 12
rect 49 8 53 10
rect 55 8 58 16
rect 60 15 65 16
rect 60 12 61 15
rect 64 12 65 15
rect 60 10 65 12
rect 69 15 74 16
rect 69 12 70 15
rect 73 12 74 15
rect 69 10 74 12
rect 60 8 64 10
<< ndc >>
rect 9 12 12 15
rect 48 12 51 15
rect 61 12 64 15
rect 70 12 73 15
<< ntransistor >>
rect 13 10 41 16
rect 44 10 46 16
rect 53 8 55 16
rect 58 8 60 16
rect 65 10 69 16
<< pdiffusion >>
rect 49 29 53 34
rect 8 27 13 29
rect 8 24 9 27
rect 12 24 13 27
rect 8 23 13 24
rect 27 23 44 29
rect 46 27 53 29
rect 46 24 48 27
rect 51 24 53 27
rect 46 23 53 24
rect 55 23 58 34
rect 60 33 64 34
rect 60 27 65 33
rect 60 24 61 27
rect 64 24 65 27
rect 60 23 65 24
rect 69 27 74 33
rect 69 24 70 27
rect 73 24 74 27
rect 69 23 74 24
<< pdc >>
rect 9 24 12 27
rect 48 24 51 27
rect 61 24 64 27
rect 70 24 73 27
<< ptransistor >>
rect 13 23 27 29
rect 44 23 46 29
rect 53 23 55 34
rect 58 23 60 34
rect 65 23 69 33
<< polysilicon >>
rect 8 43 60 45
rect 8 40 13 43
rect 8 37 9 40
rect 12 37 13 40
rect 36 39 55 40
rect 24 38 29 39
rect 8 36 13 37
rect 16 36 21 37
rect 16 33 17 36
rect 20 33 21 36
rect 24 35 25 38
rect 28 36 29 38
rect 36 36 37 39
rect 40 38 55 39
rect 40 36 41 38
rect 51 36 55 38
rect 28 35 32 36
rect 36 35 41 36
rect 24 34 32 35
rect 53 34 55 36
rect 58 34 60 43
rect 16 31 21 33
rect 30 32 32 34
rect 13 29 27 31
rect 30 30 46 32
rect 44 29 46 30
rect 65 33 69 35
rect 13 21 27 23
rect 13 16 41 18
rect 44 16 46 23
rect 53 16 55 23
rect 58 16 60 23
rect 65 21 69 23
rect 77 21 82 22
rect 65 18 78 21
rect 81 18 82 21
rect 65 16 69 18
rect 77 17 82 18
rect 13 8 41 10
rect 44 8 46 10
rect 65 8 69 10
rect 20 6 25 8
rect 30 7 35 8
rect 53 6 55 8
rect 58 6 60 8
rect 20 3 21 6
rect 24 3 25 6
rect 20 2 25 3
<< pc >>
rect 9 37 12 40
rect 17 33 20 36
rect 25 35 28 38
rect 37 36 40 39
rect 78 18 81 21
rect 21 3 24 6
<< m1 >>
rect 9 40 12 41
rect 8 37 9 40
rect 32 39 36 40
rect 56 39 60 40
rect 24 38 29 39
rect 8 36 12 37
rect 16 36 21 37
rect 16 33 17 36
rect 20 33 21 36
rect 24 35 25 38
rect 28 35 29 38
rect 32 36 37 39
rect 40 36 41 39
rect 56 36 57 39
rect 24 34 29 35
rect 16 32 21 33
rect 26 33 29 34
rect 79 35 84 40
rect 26 30 73 33
rect 79 32 80 35
rect 83 32 84 35
rect 69 28 73 30
rect 69 27 74 28
rect 8 24 9 27
rect 12 24 13 27
rect 47 24 48 27
rect 51 24 52 27
rect 60 24 61 27
rect 64 24 65 27
rect 69 24 70 27
rect 73 24 74 27
rect 9 22 13 24
rect 9 19 24 22
rect 9 15 12 16
rect 8 12 9 15
rect 12 12 13 15
rect 8 11 13 12
rect 8 5 9 8
rect 8 4 12 5
rect 21 6 24 19
rect 48 15 51 24
rect 69 23 74 24
rect 70 16 73 23
rect 78 21 81 22
rect 60 15 65 16
rect 60 12 61 15
rect 64 12 65 15
rect 69 15 74 16
rect 69 12 70 15
rect 73 12 74 15
rect 48 10 51 12
rect 78 8 81 18
rect 21 2 24 3
<< m2c >>
rect 17 33 20 36
rect 57 36 60 39
rect 80 32 83 35
rect 9 24 12 27
rect 61 24 64 27
rect 9 12 12 15
rect 9 5 12 8
rect 61 12 64 15
rect 48 7 51 10
rect 78 5 81 8
<< m2 >>
rect 56 39 61 40
rect 16 36 21 37
rect 16 33 17 36
rect 20 33 21 36
rect 56 36 57 39
rect 60 36 61 39
rect 56 35 61 36
rect 79 35 84 40
rect 16 32 21 33
rect 4 30 18 32
rect 4 15 6 30
rect 57 28 59 35
rect 79 32 80 35
rect 83 32 84 35
rect 79 31 84 32
rect 8 27 13 28
rect 57 27 65 28
rect 8 24 9 27
rect 12 24 61 27
rect 64 24 65 27
rect 8 23 13 24
rect 60 23 65 24
rect 8 15 65 16
rect 80 15 83 31
rect 4 13 9 15
rect 8 12 9 13
rect 12 14 61 15
rect 12 12 13 14
rect 8 11 13 12
rect 60 12 61 14
rect 64 12 83 15
rect 60 11 65 12
rect 47 10 52 11
rect 47 9 48 10
rect 8 8 48 9
rect 8 5 9 8
rect 12 7 48 8
rect 51 9 52 10
rect 51 8 82 9
rect 51 7 78 8
rect 12 5 13 7
rect 47 6 52 7
rect 8 4 13 5
rect 77 5 78 7
rect 81 5 82 8
rect 77 4 82 5
<< labels >>
rlabel space 0 0 88 48 6 prboundary
rlabel polysilicon 78 22 78 22 3 out
rlabel polysilicon 78 18 78 18 3 out
rlabel polysilicon 82 19 82 19 3 out
rlabel polysilicon 59 35 59 35 3 in(0)
rlabel polysilicon 41 39 41 39 3 in(1)
rlabel polysilicon 66 9 66 9 3 out
rlabel ndiffusion 70 11 70 11 3 #7
rlabel polysilicon 66 17 66 17 3 out
rlabel polysilicon 66 19 66 19 3 out
rlabel polysilicon 66 22 66 22 3 out
rlabel polysilicon 54 35 54 35 3 in(1)
rlabel ntransistor 66 11 66 11 3 out
rlabel polysilicon 66 34 66 34 3 out
rlabel polysilicon 52 37 52 37 3 in(1)
rlabel polysilicon 37 36 37 36 3 in(1)
rlabel polysilicon 37 37 37 37 3 in(1)
rlabel ndiffusion 61 9 61 9 3 GND
rlabel ndiffusion 61 11 61 11 3 GND
rlabel polysilicon 59 17 59 17 3 in(0)
rlabel ptransistor 66 24 66 24 3 out
rlabel pdiffusion 50 30 50 30 3 out
rlabel ntransistor 59 9 59 9 3 in(0)
rlabel pdiffusion 61 28 61 28 3 Vdd
rlabel pdiffusion 61 34 61 34 3 Vdd
rlabel polysilicon 29 37 29 37 3 #7
rlabel polysilicon 54 17 54 17 3 in(1)
rlabel ptransistor 59 24 59 24 3 in(0)
rlabel polysilicon 45 30 45 30 3 #7
rlabel polysilicon 59 7 59 7 3 in(0)
rlabel ntransistor 54 9 54 9 3 in(1)
rlabel ndiffusion 52 13 52 13 3 out
rlabel polysilicon 37 40 37 40 3 in(1)
rlabel ndiffusion 50 9 50 9 3 out
rlabel ptransistor 54 24 54 24 3 in(1)
rlabel polysilicon 54 7 54 7 3 in(1)
rlabel polysilicon 25 4 25 4 3 Vdd
rlabel polysilicon 31 8 31 8 3 Vdd
rlabel ndiffusion 47 11 47 11 3 out
rlabel ndiffusion 47 13 47 13 3 out
rlabel ndiffusion 47 16 47 16 3 out
rlabel pdiffusion 47 24 47 24 3 out
rlabel pdiffusion 47 25 47 25 3 out
rlabel pdiffusion 47 28 47 28 3 out
rlabel polysilicon 31 31 31 31 3 #7
rlabel polysilicon 31 33 31 33 3 #7
rlabel polysilicon 45 9 45 9 3 #7
rlabel ntransistor 45 11 45 11 3 #7
rlabel polysilicon 45 17 45 17 3 #7
rlabel ptransistor 45 24 45 24 3 #7
rlabel polysilicon 21 3 21 3 3 Vdd
rlabel polysilicon 21 4 21 4 3 Vdd
rlabel polysilicon 21 7 21 7 3 Vdd
rlabel polysilicon 17 32 17 32 3 GND
rlabel polysilicon 13 38 13 38 3 in(0)
rlabel polysilicon 14 9 14 9 3 Vdd
rlabel ntransistor 14 11 14 11 3 Vdd
rlabel polysilicon 14 17 14 17 3 Vdd
rlabel polysilicon 14 22 14 22 3 GND
rlabel ptransistor 14 24 14 24 3 GND
rlabel polysilicon 14 30 14 30 3 GND
rlabel ndiffusion 9 11 9 11 3 GND
rlabel polysilicon 9 41 9 41 3 in(0)
rlabel polysilicon 9 44 9 44 3 in(0)
rlabel m1 74 13 74 13 3 #7
rlabel m1 74 25 74 25 3 #7
rlabel ndc 71 13 71 13 3 #7
rlabel pdc 71 25 71 25 3 #7
rlabel m1 41 37 41 37 3 in(1)
port 1 e
rlabel m1 70 13 70 13 3 #7
rlabel pc 79 19 79 19 3 out
port 2 e
rlabel m1 79 22 79 22 3 out
port 2 e
rlabel m1 70 25 70 25 3 #7
rlabel m1 70 28 70 28 3 #7
rlabel m1 70 29 70 29 3 #7
rlabel pc 38 37 38 37 3 in(1)
port 1 e
rlabel m1 71 17 71 17 3 #7
rlabel m1 33 37 33 37 3 in(1)
port 1 e
rlabel m1 70 16 70 16 3 #7
rlabel m1 70 24 70 24 3 #7
rlabel m1 27 34 27 34 3 #7
rlabel m1 29 36 29 36 3 #7
rlabel m1 61 16 61 16 3 GND
rlabel m1 61 25 61 25 3 Vdd
rlabel pc 26 36 26 36 3 #7
rlabel m1 25 35 25 35 3 #7
rlabel m1 25 36 25 36 3 #7
rlabel m1 33 40 33 40 3 in(1)
port 1 e
rlabel m1 52 25 52 25 3 out
port 2 e
rlabel m1 79 9 79 9 3 out
port 2 e
rlabel ndc 49 13 49 13 3 out
port 2 e
rlabel m1 49 16 49 16 3 out
port 2 e
rlabel pdc 49 25 49 25 3 out
port 2 e
rlabel m1 25 39 25 39 3 #7
rlabel m1 48 25 48 25 3 out
port 2 e
rlabel m1 49 11 49 11 3 out
port 2 e
rlabel m1 27 31 27 31 3 #7
rlabel m1 22 3 22 3 3 Vdd
rlabel pc 22 4 22 4 3 Vdd
rlabel m1 22 7 22 7 3 Vdd
rlabel m1 10 16 10 16 3 GND
rlabel m1 10 20 10 20 3 Vdd
rlabel m1 10 23 10 23 3 Vdd
rlabel pc 10 38 10 38 3 in(0)
port 3 e
rlabel m1 10 41 10 41 3 in(0)
port 3 e
rlabel m1 9 37 9 37 3 in(0)
port 3 e
rlabel m1 9 38 9 38 3 in(0)
port 3 e
rlabel m2 84 33 84 33 3 GND
rlabel m2c 81 33 81 33 3 GND
rlabel m2 65 13 65 13 3 GND
rlabel m2 80 32 80 32 3 GND
rlabel m2 80 33 80 33 3 GND
rlabel m2 82 6 82 6 3 out
port 2 e
rlabel m2c 62 13 62 13 3 GND
rlabel m2 61 24 61 24 3 Vdd
rlabel m2 80 36 80 36 3 GND
rlabel m2c 79 6 79 6 3 out
port 2 e
rlabel m2 61 12 61 12 3 GND
rlabel m2 61 13 61 13 3 GND
rlabel m2 58 28 58 28 3 Vdd
rlabel m2 58 29 58 29 3 Vdd
rlabel m2 78 5 78 5 3 out
port 2 e
rlabel m2 78 6 78 6 3 out
port 2 e
rlabel m2 57 36 57 36 3 Vdd
rlabel m2 61 37 61 37 3 Vdd
rlabel m2 65 25 65 25 3 Vdd
rlabel m2c 58 37 58 37 3 Vdd
rlabel m2 52 8 52 8 3 out
port 2 e
rlabel m2 52 9 52 9 3 out
port 2 e
rlabel m2 52 10 52 10 3 out
port 2 e
rlabel m2 48 10 48 10 3 out
port 2 e
rlabel m2 48 11 48 11 3 out
port 2 e
rlabel m2c 62 25 62 25 3 Vdd
rlabel m2 21 34 21 34 3 GND
rlabel m2 57 37 57 37 3 Vdd
rlabel m2 57 40 57 40 3 Vdd
rlabel m2 48 7 48 7 3 out
port 2 e
rlabel m2c 49 8 49 8 3 out
port 2 e
rlabel m2 81 16 81 16 3 GND
rlabel m2 13 25 13 25 3 Vdd
rlabel m2c 18 34 18 34 3 GND
rlabel m2 13 6 13 6 3 out
port 2 e
rlabel m2 13 8 13 8 3 out
port 2 e
rlabel m2 13 13 13 13 3 GND
rlabel m2 13 15 13 15 3 GND
rlabel m2c 10 25 10 25 3 Vdd
rlabel m2 17 33 17 33 3 GND
rlabel m2 17 34 17 34 3 GND
rlabel m2 17 37 17 37 3 GND
rlabel m2c 10 6 10 6 3 out
port 2 e
rlabel m2c 10 13 10 13 3 GND
rlabel m2 9 16 9 16 3 GND
rlabel m2 9 24 9 24 3 Vdd
rlabel m2 9 25 9 25 3 Vdd
rlabel m2 9 28 9 28 3 Vdd
rlabel m2 9 5 9 5 3 out
port 2 e
rlabel m2 9 6 9 6 3 out
port 2 e
rlabel m2 9 9 9 9 3 out
port 2 e
rlabel m2 9 12 9 12 3 GND
rlabel m2 9 13 9 13 3 GND
rlabel m2 5 14 5 14 3 GND
rlabel m2 5 16 5 16 3 GND
rlabel m2 5 31 5 31 3 GND
<< end >>
