magic
tech sky130l
timestamp 1734214594
<< ndiffusion >>
rect 8 15 13 24
rect 8 12 9 15
rect 12 12 13 15
rect 8 4 13 12
rect 15 4 20 24
rect 22 8 27 24
rect 22 5 23 8
rect 26 5 27 8
rect 22 4 27 5
<< ndc >>
rect 9 12 12 15
rect 23 5 26 8
<< ntransistor >>
rect 13 4 15 24
rect 20 4 22 24
<< pdiffusion >>
rect 8 35 13 46
rect 8 32 9 35
rect 12 32 13 35
rect 8 31 13 32
rect 15 42 20 46
rect 15 39 16 42
rect 19 39 20 42
rect 15 31 20 39
rect 22 35 27 46
rect 22 32 23 35
rect 26 32 27 35
rect 22 31 27 32
<< pdc >>
rect 9 32 12 35
rect 16 39 19 42
rect 23 32 26 35
<< ptransistor >>
rect 13 31 15 46
rect 20 31 22 46
<< polysilicon >>
rect 32 60 37 61
rect 32 57 33 60
rect 36 57 37 60
rect 32 56 37 57
rect 8 53 13 54
rect 8 50 9 53
rect 12 51 13 53
rect 12 50 15 51
rect 32 50 34 56
rect 8 49 15 50
rect 13 46 15 49
rect 20 48 34 50
rect 20 46 22 48
rect 13 24 15 31
rect 20 24 22 31
rect 13 2 15 4
rect 20 2 22 4
<< pc >>
rect 33 57 36 60
rect 9 50 12 53
<< m1 >>
rect 33 61 37 65
rect 6 54 13 61
rect 20 60 27 61
rect 20 57 22 60
rect 25 57 27 60
rect 20 56 27 57
rect 31 60 39 61
rect 31 57 33 60
rect 36 57 39 60
rect 6 53 12 54
rect 6 50 9 53
rect 6 48 12 50
rect 16 53 26 56
rect 16 42 19 53
rect 31 50 39 57
rect 15 39 16 42
rect 19 39 20 42
rect 8 32 9 35
rect 12 32 23 35
rect 26 32 27 35
rect 9 15 12 32
rect 9 8 12 12
rect 6 2 12 8
rect 22 5 23 8
rect 26 5 32 8
rect 35 5 36 8
rect 30 2 36 5
<< m2c >>
rect 22 57 25 60
rect 32 5 35 8
<< m2 >>
rect 20 60 27 61
rect 20 57 22 60
rect 25 57 27 60
rect 20 56 27 57
rect 30 8 36 16
rect 30 5 32 8
rect 35 5 36 8
rect 30 2 36 5
<< labels >>
rlabel polysilicon 33 51 33 51 3 B
rlabel polysilicon 33 57 33 57 3 B
rlabel polysilicon 33 58 33 58 3 B
rlabel polysilicon 33 61 33 61 3 B
rlabel pdiffusion 23 32 23 32 3 Y
rlabel pdiffusion 23 33 23 33 3 Y
rlabel pdiffusion 23 36 23 36 3 Y
rlabel polysilicon 21 3 21 3 3 B
rlabel ntransistor 21 5 21 5 3 B
rlabel polysilicon 21 25 21 25 3 B
rlabel ptransistor 21 32 21 32 3 B
rlabel polysilicon 21 47 21 47 3 B
rlabel polysilicon 21 49 21 49 3 B
rlabel ndiffusion 13 13 13 13 3 Y
rlabel polysilicon 13 51 13 51 3 A
rlabel polysilicon 13 52 13 52 3 A
rlabel polysilicon 14 3 14 3 3 A
rlabel ntransistor 14 5 14 5 3 A
rlabel polysilicon 14 25 14 25 3 A
rlabel ptransistor 14 32 14 32 3 A
rlabel polysilicon 14 47 14 47 3 A
rlabel ndiffusion 9 5 9 5 3 Y
rlabel ndiffusion 9 13 9 13 3 Y
rlabel ndiffusion 9 16 9 16 3 Y
rlabel pdiffusion 9 32 9 32 3 Y
rlabel pdiffusion 9 36 9 36 3 Y
rlabel polysilicon 9 50 9 50 3 A
rlabel polysilicon 9 51 9 51 3 A
rlabel polysilicon 9 54 9 54 3 A
rlabel m1 37 58 37 58 3 B
port 1 e
rlabel pc 34 58 34 58 3 B
port 1 e
rlabel m1 32 51 32 51 3 B
port 1 e
rlabel m1 32 58 32 58 3 B
port 1 e
rlabel m1 34 62 34 62 3 B
port 1 e
rlabel m1 32 61 32 61 3 B
port 1 e
rlabel m1 27 33 27 33 3 Y
port 2 e
rlabel pdc 24 33 24 33 3 Y
port 2 e
rlabel m1 13 33 13 33 3 Y
port 2 e
rlabel m1 10 9 10 9 3 Y
port 2 e
rlabel ndc 10 13 10 13 3 Y
port 2 e
rlabel m1 10 16 10 16 3 Y
port 2 e
rlabel pdc 10 33 10 33 3 Y
port 2 e
rlabel m1 9 33 9 33 3 Y
port 2 e
rlabel pc 10 51 10 51 3 A
port 3 e
rlabel m1 7 3 7 3 3 Y
port 2 e
rlabel m1 7 49 7 49 3 A
port 3 e
rlabel m1 7 51 7 51 3 A
port 3 e
rlabel m1 7 54 7 54 3 A
port 3 e
rlabel m1 7 55 7 55 3 A
port 3 e
rlabel m2 36 6 36 6 3 GND
rlabel m2c 33 6 33 6 3 GND
rlabel m2 31 3 31 3 3 GND
rlabel m2 31 6 31 6 3 GND
rlabel m2 31 9 31 9 3 GND
rlabel m2 26 58 26 58 3 Vdd
rlabel m2c 23 58 23 58 3 Vdd
rlabel m2 21 57 21 57 3 Vdd
rlabel m2 21 58 21 58 3 Vdd
rlabel m2 21 61 21 61 3 Vdd
<< end >>
