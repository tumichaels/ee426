magic
tech sky130l
timestamp 1731038682
<< ndiffusion >>
rect 8 11 13 12
rect 8 7 9 11
rect 12 7 13 11
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
rect 22 11 27 12
rect 22 7 23 11
rect 26 7 27 11
rect 22 6 27 7
<< ndc >>
rect 9 7 12 11
rect 16 8 19 11
rect 23 7 26 11
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
<< pdiffusion >>
rect 8 33 13 34
rect 8 30 9 33
rect 12 30 13 33
rect 8 19 13 30
rect 15 19 20 34
rect 22 25 27 34
rect 22 22 23 25
rect 26 22 27 25
rect 22 19 27 22
<< pdc >>
rect 9 30 12 33
rect 23 22 26 25
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
<< polysilicon >>
rect 8 42 13 43
rect 23 42 28 43
rect 8 39 9 42
rect 12 39 15 42
rect 8 38 15 39
rect 13 34 15 38
rect 20 39 24 42
rect 27 39 28 42
rect 20 38 28 39
rect 20 34 22 38
rect 13 12 15 19
rect 20 12 22 19
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 9 39 12 42
rect 24 39 27 42
<< m1 >>
rect 8 43 12 48
rect 16 47 20 48
rect 16 44 17 47
rect 16 43 20 44
rect 8 42 13 43
rect 8 39 9 42
rect 12 39 13 42
rect 8 38 13 39
rect 8 33 13 34
rect 8 30 9 33
rect 12 32 13 33
rect 16 32 19 43
rect 23 42 28 43
rect 32 42 36 48
rect 23 39 24 42
rect 27 39 35 42
rect 23 38 28 39
rect 12 30 19 32
rect 8 29 19 30
rect 23 25 27 27
rect 26 22 27 25
rect 23 19 27 22
rect 15 15 36 19
rect 8 11 12 12
rect 8 7 9 11
rect 15 11 20 15
rect 15 8 16 11
rect 19 8 20 11
rect 15 7 20 8
rect 23 11 27 12
rect 26 7 27 11
rect 8 4 12 7
rect 23 4 27 7
rect 8 1 9 4
rect 12 1 27 4
rect 8 0 27 1
rect 32 0 36 15
<< m2c >>
rect 17 44 20 47
rect 9 1 12 4
<< m2 >>
rect 16 47 21 48
rect 16 44 17 47
rect 20 44 21 47
rect 16 43 21 44
rect 8 4 13 5
rect 8 1 9 4
rect 12 1 13 4
rect 8 0 13 1
<< labels >>
rlabel ndiffusion 23 7 23 7 3 GND
rlabel pdiffusion 23 20 23 20 3 Y
rlabel polysilicon 21 13 21 13 3 B
rlabel polysilicon 21 18 21 18 3 B
rlabel ndiffusion 16 7 16 7 3 Y
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 17 45 17 45 3 Vdd
port 3 e
rlabel m1 9 45 9 45 3 A
port 5 e
rlabel m1 9 1 9 1 3 GND
port 4 e
rlabel m1 33 1 33 1 3 Y
port 1 e
rlabel m1 33 45 33 45 3 B
port 2 e
<< end >>
