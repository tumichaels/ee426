magic
tech sky130l
timestamp 1731029939
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 23 13 27
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 26 20 27
rect 15 23 16 26
rect 19 23 20 26
rect 15 19 20 23
<< pdc >>
rect 9 20 12 23
rect 16 23 19 26
<< ptransistor >>
rect 13 19 15 27
<< polysilicon >>
rect 13 27 15 29
rect 13 17 15 19
rect 23 17 28 18
rect 13 15 24 17
rect 13 12 15 15
rect 23 14 24 15
rect 27 14 28 17
rect 23 13 28 14
rect 13 4 15 6
<< pc >>
rect 24 14 27 17
<< m1 >>
rect 7 31 12 32
rect 7 28 9 31
rect 7 27 12 28
rect 16 31 28 32
rect 16 28 24 31
rect 27 28 28 31
rect 16 26 19 28
rect 9 23 12 24
rect 16 22 19 23
rect 9 10 12 20
rect 19 14 24 17
rect 27 14 28 17
rect 7 7 9 9
rect 7 4 12 7
rect 16 10 19 11
rect 19 8 28 10
rect 19 7 24 8
rect 16 6 19 7
rect 23 5 24 7
rect 27 5 28 8
rect 23 4 28 5
<< m2c >>
rect 9 28 12 31
rect 24 28 27 31
rect 16 14 19 17
rect 24 5 27 8
<< m2 >>
rect 8 31 13 32
rect 8 28 9 31
rect 12 28 13 31
rect 8 27 13 28
rect 23 31 28 32
rect 23 28 24 31
rect 27 28 28 31
rect 23 27 28 28
rect 9 17 11 27
rect 15 17 20 18
rect 9 15 16 17
rect 15 14 16 15
rect 19 14 20 17
rect 15 13 20 14
rect 23 8 28 9
rect 23 5 24 8
rect 27 5 28 8
rect 23 4 28 5
<< labels >>
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel m1 17 29 17 29 3 Vdd
port 2 e
rlabel m1 9 5 9 5 3 Y
port 3 e
rlabel m1 9 29 9 29 3 A
port 4 e
rlabel m1 7 28 9 32 4 A
rlabel m2 26 5 26 5 8 GND
<< end >>
