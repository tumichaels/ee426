magic
tech sky130l
timestamp 1731040963
<< ndiffusion >>
rect 8 11 13 12
rect 8 8 9 11
rect 12 8 13 11
rect 8 6 13 8
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 8 12 11
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 23 13 25
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 24 20 25
rect 15 21 16 24
rect 19 21 20 24
rect 15 19 20 21
<< pdc >>
rect 9 20 12 23
rect 16 21 19 24
<< ptransistor >>
rect 13 19 15 25
<< polysilicon >>
rect 13 25 15 27
rect 13 17 15 19
rect 23 18 28 19
rect 23 17 24 18
rect 13 15 24 17
rect 27 15 28 18
rect 13 12 15 15
rect 23 14 28 15
rect 13 4 15 6
<< pc >>
rect 24 15 27 18
<< m1 >>
rect 7 31 12 32
rect 7 28 9 31
rect 16 28 22 31
rect 16 24 19 28
rect 9 23 12 24
rect 15 21 16 24
rect 19 21 20 24
rect 9 11 12 20
rect 23 18 28 19
rect 19 15 24 18
rect 27 15 28 18
rect 23 14 28 15
rect 15 8 16 11
rect 19 8 28 11
rect 7 4 12 8
rect 27 5 28 8
rect 24 4 28 5
<< m2c >>
rect 9 28 12 31
rect 22 28 25 31
rect 16 15 19 18
rect 24 5 27 8
<< m2 >>
rect 8 31 13 32
rect 8 28 9 31
rect 12 28 13 31
rect 8 27 13 28
rect 21 31 26 32
rect 21 28 22 31
rect 25 28 26 31
rect 21 27 26 28
rect 9 18 12 27
rect 15 18 20 19
rect 9 15 16 18
rect 19 15 20 18
rect 15 14 20 15
rect 23 8 28 9
rect 23 5 24 8
rect 27 5 28 8
rect 23 4 28 5
<< labels >>
rlabel space 0 0 32 36 6 prboundary
rlabel polysilicon 24 18 24 18 3 in(0)
rlabel ndiffusion 16 7 16 7 3 GND
rlabel ndiffusion 16 12 16 12 3 GND
rlabel ndiffusion 13 9 13 9 3 out
rlabel pdiffusion 16 20 16 20 3 Vdd
rlabel pdiffusion 16 25 16 25 3 Vdd
rlabel pdiffusion 13 21 13 21 3 out
rlabel polysilicon 14 5 14 5 3 in(0)
rlabel ntransistor 14 7 14 7 3 in(0)
rlabel polysilicon 14 13 14 13 3 in(0)
rlabel polysilicon 14 16 14 16 3 in(0)
rlabel polysilicon 14 18 14 18 3 in(0)
rlabel ptransistor 14 20 14 20 3 in(0)
rlabel polysilicon 14 26 14 26 3 in(0)
rlabel ndiffusion 9 7 9 7 3 out
rlabel ndiffusion 9 9 9 9 3 out
rlabel ndiffusion 9 12 9 12 3 out
rlabel pdiffusion 9 20 9 20 3 out
rlabel pdiffusion 9 21 9 21 3 out
rlabel pdiffusion 9 24 9 24 3 out
rlabel m1 28 16 28 16 3 in(0)
port 1 e
rlabel m1 24 15 24 15 3 in(0)
port 1 e
rlabel pc 25 16 25 16 3 in(0)
port 1 e
rlabel m1 24 19 24 19 3 in(0)
port 1 e
rlabel m1 20 9 20 9 3 GND
rlabel m1 20 22 20 22 3 Vdd
rlabel ndc 17 9 17 9 3 GND
rlabel pdc 17 22 17 22 3 Vdd
rlabel m1 17 25 17 25 3 Vdd
rlabel m1 17 29 17 29 3 Vdd
rlabel m1 16 9 16 9 3 GND
rlabel m1 16 22 16 22 3 Vdd
rlabel m1 25 5 25 5 3 GND
rlabel ndc 10 9 10 9 3 out
port 2 e
rlabel m1 10 12 10 12 3 out
port 2 e
rlabel pdc 10 21 10 21 3 out
port 2 e
rlabel m1 10 24 10 24 3 out
port 2 e
rlabel m1 8 5 8 5 3 out
port 2 e
rlabel m1 8 29 8 29 3 in(0)
port 1 e
rlabel m1 8 32 8 32 3 in(0)
port 1 e
rlabel m2 28 6 28 6 3 GND
rlabel m2 26 29 26 29 3 Vdd
rlabel m2c 25 6 25 6 3 GND
rlabel m2 22 28 22 28 3 Vdd
rlabel m2c 23 29 23 29 3 Vdd
rlabel m2 24 5 24 5 3 GND
rlabel m2 24 6 24 6 3 GND
rlabel m2 24 9 24 9 3 GND
rlabel m2 22 29 22 29 3 Vdd
rlabel m2 20 16 20 16 3 in(0)
port 1 e
rlabel m2 16 19 16 19 3 in(0)
port 1 e
rlabel m2 16 15 16 15 3 in(0)
port 1 e
rlabel m2c 17 16 17 16 3 in(0)
port 1 e
rlabel m2 13 29 13 29 3 in(0)
port 1 e
rlabel m2 22 32 22 32 3 Vdd
rlabel m2 10 16 10 16 3 in(0)
port 1 e
rlabel m2 10 19 10 19 3 in(0)
port 1 e
rlabel m2c 10 29 10 29 3 in(0)
port 1 e
rlabel m2 9 28 9 28 3 in(0)
port 1 e
rlabel m2 9 29 9 29 3 in(0)
port 1 e
rlabel m2 9 32 9 32 3 in(0)
port 1 e
<< end >>
