magic
tech sky130l
timestamp 1730909014
<< ndiffusion >>
rect 8 15 13 16
rect 8 11 9 15
rect 12 11 13 15
rect 8 10 13 11
rect 15 15 20 16
rect 15 12 16 15
rect 19 12 20 15
rect 15 10 20 12
rect 22 15 27 16
rect 22 11 23 15
rect 26 11 27 15
rect 22 10 27 11
<< ndc >>
rect 9 11 12 15
rect 16 12 19 15
rect 23 11 26 15
<< ntransistor >>
rect 13 10 15 16
rect 20 10 22 16
<< pdiffusion >>
rect 8 37 13 38
rect 8 34 9 37
rect 12 34 13 37
rect 8 23 13 34
rect 15 23 20 38
rect 22 29 27 38
rect 22 26 23 29
rect 26 26 27 29
rect 22 23 27 26
<< pdc >>
rect 9 34 12 37
rect 23 26 26 29
<< ptransistor >>
rect 13 23 15 38
rect 20 23 22 38
<< polysilicon >>
rect 8 46 13 47
rect 23 46 28 47
rect 8 43 9 46
rect 12 43 15 46
rect 8 42 15 43
rect 13 38 15 42
rect 20 43 24 46
rect 27 43 28 46
rect 20 42 28 43
rect 20 38 22 42
rect 13 16 15 23
rect 20 16 22 23
rect 13 8 15 10
rect 20 8 22 10
<< pc >>
rect 9 43 12 46
rect 24 43 27 46
<< m1 >>
rect 8 47 12 52
rect 8 46 13 47
rect 8 43 9 46
rect 12 43 13 46
rect 8 42 13 43
rect 8 37 13 38
rect 8 34 9 37
rect 12 36 13 37
rect 16 36 20 52
rect 24 47 28 52
rect 23 46 28 47
rect 23 43 24 46
rect 27 43 28 46
rect 23 42 28 43
rect 12 34 20 36
rect 8 33 20 34
rect 23 29 27 31
rect 26 26 27 29
rect 23 23 27 26
rect 32 23 36 52
rect 15 19 36 23
rect 8 15 12 16
rect 8 11 9 15
rect 15 15 20 19
rect 15 12 16 15
rect 19 12 20 15
rect 15 11 20 12
rect 23 15 27 16
rect 26 11 27 15
rect 8 8 12 11
rect 23 8 27 11
rect 8 4 27 8
<< labels >>
rlabel space 0 0 40 56 6 prboundary
rlabel ndiffusion 23 11 23 11 3 GND
rlabel ndiffusion 23 12 23 12 3 GND
rlabel ndiffusion 23 16 23 16 3 GND
rlabel pdiffusion 23 24 23 24 3 Y
rlabel pdiffusion 23 27 23 27 3 Y
rlabel pdiffusion 23 30 23 30 3 Y
rlabel polysilicon 21 9 21 9 3 B
rlabel ntransistor 21 11 21 11 3 B
rlabel polysilicon 21 17 21 17 3 B
rlabel ptransistor 21 24 21 24 3 B
rlabel polysilicon 21 39 21 39 3 B
rlabel polysilicon 21 43 21 43 3 B
rlabel polysilicon 21 44 21 44 3 B
rlabel ndiffusion 16 11 16 11 3 Y
rlabel ndiffusion 13 12 13 12 3 GND
rlabel polysilicon 14 9 14 9 3 A
rlabel ntransistor 14 11 14 11 3 A
rlabel polysilicon 14 17 14 17 3 A
rlabel ptransistor 14 24 14 24 3 A
rlabel polysilicon 14 39 14 39 3 A
rlabel ndiffusion 9 11 9 11 3 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m1 33 24 33 24 3 Y
port 1 e
rlabel m1 28 44 28 44 3 B
port 2 e
rlabel m1 27 27 27 27 3 Y
port 1 e
rlabel pc 25 44 25 44 3 B
port 2 e
rlabel m1 25 48 25 48 3 B
port 2 e
rlabel m1 27 12 27 12 3 GND
rlabel m1 24 24 24 24 3 Y
port 1 e
rlabel pdc 24 27 24 27 3 Y
port 1 e
rlabel m1 24 30 24 30 3 Y
port 1 e
rlabel m1 24 43 24 43 3 B
port 2 e
rlabel m1 24 44 24 44 3 B
port 2 e
rlabel m1 24 47 24 47 3 B
port 2 e
rlabel ndc 24 12 24 12 3 GND
rlabel m1 20 13 20 13 3 Y
port 1 e
rlabel m1 24 16 24 16 3 GND
rlabel ndc 17 13 17 13 3 Y
port 1 e
rlabel m1 17 37 17 37 3 Vdd
rlabel m1 16 12 16 12 3 Y
port 1 e
rlabel m1 16 13 16 13 3 Y
port 1 e
rlabel m1 16 16 16 16 3 Y
port 1 e
rlabel m1 16 20 16 20 3 Y
port 1 e
rlabel m1 24 9 24 9 3 GND
rlabel m1 13 35 13 35 3 Vdd
rlabel m1 13 37 13 37 3 Vdd
rlabel m1 13 44 13 44 3 A
port 3 e
rlabel ndc 10 12 10 12 3 GND
rlabel pdc 10 35 10 35 3 Vdd
rlabel pc 10 44 10 44 3 A
port 3 e
rlabel m1 9 5 9 5 3 GND
rlabel m1 9 9 9 9 3 GND
rlabel m1 9 12 9 12 3 GND
rlabel m1 9 16 9 16 3 GND
rlabel m1 9 34 9 34 3 Vdd
rlabel m1 9 35 9 35 3 Vdd
rlabel m1 9 38 9 38 3 Vdd
rlabel m1 9 43 9 43 3 A
port 3 e
rlabel m1 9 44 9 44 3 A
port 3 e
rlabel m1 9 47 9 47 3 A
port 3 e
rlabel m1 9 48 9 48 3 A
port 3 e
<< end >>
