magic
tech TSMC180
timestamp 1734147306
<< ndiffusion >>
rect 6 9 12 12
rect 14 9 20 12
<< ntransistor >>
rect 12 9 14 12
<< pdiffusion >>
rect 6 28 12 31
rect 14 28 20 31
<< ptransistor >>
rect 12 28 14 31
<< polysilicon >>
rect 12 31 14 34
rect 12 25 14 28
rect 12 12 14 15
rect 12 6 14 9
<< m1 >>
rect 6 37 9 40
rect 24 37 27 40
<< labels >>
rlabel ndiffusion 15 10 15 10 3 Y
rlabel pdiffusion 15 29 15 29 3 x
rlabel polysilicon 13 13 13 13 3 x
rlabel polysilicon 13 26 13 26 3 x
rlabel ndiffusion 7 10 7 10 3 GND
rlabel pdiffusion 7 29 7 29 3 Vdd
rlabel m1 25 38 25 38 3 GND
port 1 e
rlabel m1 7 38 7 38 3 Vdd
port 3 e
<< end >>
