magic
tech sky130l
timestamp 1726533950
<< polysilicon >>
rect -45 104 -34 109
rect -45 88 -34 93
rect -45 51 -34 56
rect -45 35 -34 40
<< pc >>
rect -42 143 -39 146
<< m1 >>
rect -13 165 -6 174
rect -43 154 -38 163
rect -43 151 -42 154
rect -39 151 -38 154
rect -43 150 -38 151
rect -43 146 -38 147
rect -43 143 -42 146
rect -39 143 -38 146
rect -43 74 -38 143
rect -43 70 -42 74
rect -39 70 -38 74
rect -43 69 -38 70
rect -34 26 -27 133
rect -13 128 -6 129
rect -13 124 -12 128
rect -7 124 -6 128
rect -13 120 -6 124
rect -13 74 -6 75
rect -13 70 -12 74
rect -7 70 -6 74
rect -13 67 -6 70
rect 8 26 15 140
<< m2c >>
rect -42 151 -39 154
rect -42 70 -39 74
rect -12 124 -7 128
rect -12 70 -7 74
<< m2 >>
rect -43 154 -38 155
rect -43 151 -42 154
rect -39 151 -38 154
rect -43 129 -38 151
rect -43 128 -6 129
rect -43 124 -12 128
rect -7 124 -6 128
rect -43 123 -6 124
rect -43 74 -6 75
rect -43 70 -42 74
rect -39 70 -12 74
rect -7 70 -6 74
rect -43 69 -6 70
use nand2  nand2_1 ../nand
timestamp 1726527220
transform 1 0 -89 0 1 100
box 44 31 104 74
use nor2  nor2_0 ../nor
timestamp 1726527990
transform 1 0 -301 0 1 -74
box 256 151 316 194
use nor2  nor2_2
timestamp 1726527990
transform 1 0 -301 0 1 -127
box 256 151 316 194
<< labels >>
rlabel polysilicon -45 35 -34 40 7 in11
rlabel polysilicon -45 51 -34 56 7 in10
rlabel polysilicon -45 88 -34 93 7 in01
rlabel polysilicon -45 104 -34 109 7 in00
rlabel m1 -13 165 -6 174 1 out
rlabel m1 -34 26 -27 133 5 Vdd!
rlabel m1 8 65 15 80 3 GND!
<< end >>
