VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005000 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 0.600000 BY 0.300000 ;
END CoreSite

LAYER li
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.056250 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.225000 ;
   PITCH 0.600000 0.600000 ;
END li

LAYER mcon
    TYPE CUT ;
    SPACING 0.225000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END mcon

LAYER met1
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.150000 ;
   AREA 0.084375 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met1

LAYER v1
    TYPE CUT ;
    SPACING 0.075000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.075000 ;
END v1

LAYER met2
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.150000 ;
   AREA 0.073125 ;
   WIDTH 0.150000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.150000 ;
   PITCH 0.300000 0.300000 ;
END met2

LAYER v2
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.300000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v2

LAYER met3
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met3

LAYER v3
    TYPE CUT ;
    SPACING 0.150000 ;
    WIDTH 0.450000 ;
    ENCLOSURE ABOVE 0.075000 0.075000 ;
    ENCLOSURE BELOW 0.075000 0.000000 ;
END v3

LAYER met4
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.300000 ;
   AREA 0.241875 ;
   WIDTH 0.300000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.300000 ;
   PITCH 0.600000 0.600000 ;
END met4

LAYER v4
    TYPE CUT ;
    SPACING 0.450000 ;
    WIDTH 1.200000 ;
    ENCLOSURE ABOVE 0.150000 0.150000 ;
    ENCLOSURE BELOW 0.000000 0.000000 ;
END v4

LAYER met5
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 1.650000 ;
   AREA 4.005000 ;
   WIDTH 1.650000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 1.650000 ;
   PITCH 3.300000 3.300000 ;
END met5

LAYER OVERLAP
   TYPE OVERLAP ;
END OVERLAP

VIA mcon_C DEFAULT
   LAYER li ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER mcon ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END mcon_C

VIA v1_C DEFAULT
   LAYER met1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_C

VIA v2_C DEFAULT
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_C

VIA v2_Ch
   LAYER met2 ;
     RECT -0.225000 -0.150000 0.225000 0.150000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Ch

VIA v2_Cv
   LAYER met2 ;
     RECT -0.150000 -0.225000 0.150000 0.225000 ;
   LAYER v2 ;
     RECT -0.150000 -0.150000 0.150000 0.150000 ;
   LAYER met3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Cv

VIA v3_C DEFAULT
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_C

VIA v3_Ch
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Ch

VIA v3_Cv
   LAYER met3 ;
     RECT -0.300000 -0.225000 0.300000 0.225000 ;
   LAYER v3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER met4 ;
     RECT -0.300000 -0.300000 0.300000 0.300000 ;
END v3_Cv

VIA v4_C DEFAULT
   LAYER met4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER v4 ;
     RECT -0.600000 -0.600000 0.600000 0.600000 ;
   LAYER met5 ;
     RECT -0.750000 -0.750000 0.750000 0.750000 ;
END v4_C

MACRO _0_0std_0_0cells_0_0FAX1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0FAX1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 10.200000 BY 8.700000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 8.325000 2.325000 8.400000 ;
        RECT 0.600000 8.100000 2.025000 8.325000 ;
        RECT 2.025000 8.100000 2.250000 8.325000 ;
        RECT 2.250000 8.100000 2.325000 8.325000 ;
        RECT 1.950000 8.025000 2.325000 8.100000 ;
        RECT 4.950000 8.325000 5.325000 8.400000 ;
        RECT 4.950000 8.100000 5.025000 8.325000 ;
        RECT 4.950000 8.025000 5.325000 8.100000 ;
        RECT 4.950000 6.525000 5.325000 6.600000 ;
        RECT 4.950000 6.300000 5.025000 6.525000 ;
        RECT 4.950000 6.225000 5.325000 6.300000 ;
        RECT 5.025000 8.100000 5.250000 8.325000 ;
        RECT 5.025000 6.600000 5.250000 8.025000 ;
        RECT 5.025000 6.300000 5.250000 6.525000 ;
        RECT 5.250000 8.100000 5.325000 8.325000 ;
        RECT 5.250000 6.300000 5.325000 6.525000 ;
        END
        ANTENNAGATEAREA 2.182500 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 6.675000 1.500000 6.900000 ;
        RECT 0.600000 6.600000 2.850000 6.675000 ;
        RECT 1.500000 6.675000 1.725000 6.900000 ;
        RECT 1.725000 6.675000 2.850000 6.900000 ;
        RECT 1.425000 6.900000 1.800000 6.975000 ;
        RECT 2.550000 7.800000 4.425000 7.875000 ;
        RECT 2.550000 7.575000 2.625000 7.800000 ;
        RECT 2.550000 7.500000 4.425000 7.575000 ;
        RECT 2.550000 6.900000 2.850000 7.500000 ;
        RECT 2.625000 7.575000 2.850000 7.800000 ;
        RECT 2.850000 7.575000 3.975000 7.800000 ;
        RECT 3.975000 7.575000 4.200000 7.800000 ;
        RECT 4.200000 7.575000 4.425000 7.800000 ;
        RECT 6.450000 7.800000 6.825000 7.875000 ;
        RECT 6.450000 7.575000 6.525000 7.800000 ;
        RECT 6.450000 7.500000 6.825000 7.575000 ;
        RECT 6.525000 7.575000 6.750000 7.800000 ;
        RECT 6.750000 7.575000 6.825000 7.800000 ;
        END
        ANTENNAGATEAREA 2.137500 ;
    END B
    PIN C
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 5.625000 4.650000 5.700000 ;
        RECT 0.600000 5.400000 1.050000 5.625000 ;
        RECT 1.050000 5.400000 1.275000 5.625000 ;
        RECT 1.275000 5.400000 4.650000 5.625000 ;
        RECT 0.975000 5.325000 1.350000 5.400000 ;
        RECT 3.900000 7.200000 4.650000 7.275000 ;
        RECT 3.900000 6.975000 3.975000 7.200000 ;
        RECT 3.900000 6.900000 4.650000 6.975000 ;
        RECT 3.975000 6.975000 4.200000 7.200000 ;
        RECT 4.200000 6.975000 4.350000 7.200000 ;
        RECT 4.350000 6.975000 4.575000 7.200000 ;
        RECT 4.575000 6.975000 4.650000 7.200000 ;
        RECT 4.425000 5.700000 4.650000 6.900000 ;
        RECT 6.075000 7.200000 6.825000 7.275000 ;
        RECT 6.075000 6.975000 6.150000 7.200000 ;
        RECT 6.075000 6.900000 6.825000 6.975000 ;
        RECT 6.150000 6.975000 6.375000 7.200000 ;
        RECT 6.375000 6.975000 6.525000 7.200000 ;
        RECT 6.525000 6.975000 6.750000 7.200000 ;
        RECT 6.750000 6.975000 6.825000 7.200000 ;
        LAYER mcon ;
        RECT 3.975000 6.975000 4.200000 7.200000 ;
        RECT 6.525000 6.975000 6.750000 7.200000 ;
        LAYER met1 ;
        RECT 3.900000 7.200000 6.825000 7.275000 ;
        RECT 3.900000 6.975000 3.975000 7.200000 ;
        RECT 3.900000 6.900000 6.825000 6.975000 ;
        RECT 3.975000 6.975000 4.200000 7.200000 ;
        RECT 4.200000 6.975000 6.525000 7.200000 ;
        RECT 6.525000 6.975000 6.750000 7.200000 ;
        RECT 6.750000 6.975000 6.825000 7.200000 ;
        END
        ANTENNAGATEAREA 1.631250 ;
    END C
    PIN YC
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 0.600000 0.750000 8.025000 0.900000 ;
        RECT 0.600000 0.675000 8.325000 0.750000 ;
        RECT 0.600000 0.600000 8.100000 0.675000 ;
        RECT 8.025000 0.750000 8.250000 0.975000 ;
        RECT 8.250000 0.750000 8.325000 0.975000 ;
        RECT 7.950000 0.975000 8.325000 1.050000 ;
        RECT 7.950000 0.900000 8.025000 0.975000 ;
        RECT 7.800000 3.300000 8.100000 3.525000 ;
        RECT 7.800000 3.075000 8.025000 3.300000 ;
        RECT 7.800000 2.850000 8.100000 3.075000 ;
        RECT 7.800000 2.775000 8.325000 2.850000 ;
        RECT 7.800000 2.550000 8.025000 2.775000 ;
        RECT 7.800000 2.475000 8.325000 2.550000 ;
        RECT 7.800000 2.250000 8.100000 2.475000 ;
        RECT 8.025000 3.075000 8.100000 3.300000 ;
        RECT 8.025000 2.550000 8.250000 2.775000 ;
        RECT 7.800000 1.950000 8.100000 2.025000 ;
        RECT 8.250000 2.550000 8.325000 2.775000 ;
        RECT 7.800000 2.025000 8.025000 2.250000 ;
        RECT 8.025000 2.025000 8.100000 2.250000 ;
        LAYER mcon ;
        RECT 8.025000 0.750000 8.250000 0.975000 ;
        RECT 8.025000 2.550000 8.250000 2.775000 ;
        LAYER met1 ;
        RECT 7.950000 0.975000 8.325000 1.050000 ;
        RECT 7.950000 0.750000 8.025000 0.975000 ;
        RECT 7.950000 0.675000 8.325000 0.750000 ;
        RECT 8.025000 1.050000 8.250000 2.475000 ;
        RECT 8.025000 0.750000 8.250000 0.975000 ;
        RECT 7.950000 2.775000 8.325000 2.850000 ;
        RECT 7.950000 2.550000 8.025000 2.775000 ;
        RECT 7.950000 2.475000 8.325000 2.550000 ;
        RECT 8.250000 0.750000 8.325000 0.975000 ;
        RECT 8.025000 2.550000 8.250000 2.775000 ;
        RECT 8.250000 2.550000 8.325000 2.775000 ;
        END
        ANTENNADIFFAREA 0.393750 ;
    END YC
    PIN YS
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER li ;
        RECT 9.375000 0.300000 9.675000 1.950000 ;
        RECT 8.550000 3.300000 8.925000 3.525000 ;
        RECT 8.550000 2.850000 8.925000 3.075000 ;
        RECT 8.550000 2.475000 9.675000 2.700000 ;
        RECT 8.550000 3.075000 8.625000 3.300000 ;
        RECT 9.075000 1.950000 9.675000 2.025000 ;
        RECT 8.625000 3.075000 8.850000 3.300000 ;
        RECT 8.550000 2.700000 9.450000 2.850000 ;
        RECT 8.850000 3.075000 8.925000 3.300000 ;
        RECT 9.075000 2.025000 9.150000 2.250000 ;
        RECT 9.150000 2.025000 9.375000 2.250000 ;
        RECT 9.075000 2.250000 9.675000 2.475000 ;
        RECT 9.375000 2.025000 9.675000 2.250000 ;
        END
        ANTENNADIFFAREA 0.393750 ;
    END YS
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 0.600000 4.575000 0.900000 4.650000 ;
        RECT 0.600000 4.350000 0.675000 4.575000 ;
        RECT 0.600000 3.750000 0.825000 4.350000 ;
        RECT 0.600000 3.675000 5.025000 3.750000 ;
        RECT 0.600000 3.450000 0.675000 3.675000 ;
        RECT 0.600000 3.375000 0.975000 3.450000 ;
        RECT 0.675000 4.350000 0.900000 4.575000 ;
        RECT 0.675000 3.450000 0.900000 3.675000 ;
        RECT 0.900000 3.525000 3.525000 3.675000 ;
        RECT 0.900000 3.450000 0.975000 3.525000 ;
        RECT 3.450000 3.450000 3.525000 3.525000 ;
        RECT 3.450000 3.375000 3.825000 3.450000 ;
        RECT 3.525000 3.450000 3.750000 3.675000 ;
        RECT 3.750000 3.525000 4.125000 3.675000 ;
        RECT 3.750000 3.450000 3.825000 3.525000 ;
        RECT 4.050000 3.450000 4.125000 3.525000 ;
        RECT 4.050000 3.375000 4.425000 3.450000 ;
        RECT 4.125000 3.450000 4.350000 3.675000 ;
        RECT 7.200000 3.000000 7.275000 3.225000 ;
        RECT 7.200000 2.925000 7.500000 3.000000 ;
        RECT 4.350000 3.525000 4.725000 3.675000 ;
        RECT 4.350000 3.450000 4.425000 3.525000 ;
        RECT 7.275000 3.000000 7.500000 3.225000 ;
        RECT 4.650000 3.450000 4.725000 3.525000 ;
        RECT 4.650000 3.375000 5.025000 3.450000 ;
        RECT 4.725000 3.450000 4.950000 3.675000 ;
        RECT 4.950000 3.450000 5.025000 3.675000 ;
        RECT 7.125000 3.675000 7.500000 3.750000 ;
        RECT 7.125000 3.450000 7.200000 3.675000 ;
        RECT 7.125000 3.375000 7.500000 3.450000 ;
        RECT 7.200000 3.450000 7.425000 3.675000 ;
        RECT 7.200000 3.225000 7.500000 3.375000 ;
        RECT 7.425000 3.450000 7.500000 3.675000 ;
        LAYER mcon ;
        RECT 0.675000 4.350000 0.900000 4.575000 ;
        RECT 4.125000 3.450000 4.350000 3.675000 ;
        RECT 7.200000 3.450000 7.425000 3.675000 ;
        LAYER met1 ;
        RECT 0.600000 4.575000 0.975000 4.650000 ;
        RECT 0.600000 4.350000 0.675000 4.575000 ;
        RECT 0.600000 4.275000 0.975000 4.350000 ;
        RECT 0.675000 4.350000 0.900000 4.575000 ;
        RECT 0.900000 4.350000 0.975000 4.575000 ;
        RECT 4.050000 3.675000 7.575000 3.750000 ;
        RECT 4.050000 3.450000 4.125000 3.675000 ;
        RECT 4.050000 3.375000 4.425000 3.450000 ;
        RECT 4.125000 3.450000 4.350000 3.675000 ;
        RECT 4.350000 3.525000 7.200000 3.675000 ;
        RECT 4.350000 3.450000 4.425000 3.525000 ;
        RECT 7.125000 3.450000 7.200000 3.525000 ;
        RECT 7.200000 3.450000 7.425000 3.675000 ;
        RECT 7.425000 3.525000 7.575000 3.675000 ;
        RECT 7.425000 3.450000 7.500000 3.525000 ;
        RECT 7.125000 3.375000 7.500000 3.450000 ;
        END
        ANTENNADIFFAREA 4.365000 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 0.600000 1.425000 0.675000 1.650000 ;
        RECT 0.600000 1.350000 3.150000 1.425000 ;
        RECT 0.675000 1.425000 0.900000 1.650000 ;
        RECT 0.900000 1.425000 3.150000 1.650000 ;
        RECT 2.325000 1.950000 2.400000 2.175000 ;
        RECT 2.325000 1.875000 2.700000 1.950000 ;
        RECT 2.400000 1.950000 2.625000 2.175000 ;
        RECT 2.625000 1.950000 3.525000 2.175000 ;
        RECT 2.925000 1.650000 3.150000 1.950000 ;
        RECT 3.525000 1.950000 3.750000 2.175000 ;
        RECT 2.325000 2.175000 2.700000 2.250000 ;
        RECT 3.750000 1.950000 4.725000 2.175000 ;
        RECT 3.450000 1.875000 3.825000 1.950000 ;
        RECT 4.725000 1.950000 4.950000 2.175000 ;
        RECT 3.450000 2.175000 3.825000 2.250000 ;
        RECT 4.950000 1.950000 5.325000 2.175000 ;
        RECT 4.650000 1.875000 5.025000 1.950000 ;
        RECT 5.325000 1.950000 5.550000 2.175000 ;
        RECT 5.550000 1.950000 5.625000 2.175000 ;
        RECT 5.250000 1.875000 5.625000 1.950000 ;
        RECT 6.900000 2.250000 7.575000 2.325000 ;
        RECT 6.900000 2.025000 6.975000 2.250000 ;
        RECT 6.900000 1.950000 7.575000 2.025000 ;
        RECT 4.650000 2.175000 5.025000 2.250000 ;
        RECT 6.975000 2.025000 7.200000 2.250000 ;
        RECT 7.200000 2.025000 7.275000 2.250000 ;
        RECT 5.250000 2.175000 5.625000 2.250000 ;
        RECT 7.275000 2.025000 7.500000 2.250000 ;
        RECT 7.500000 2.025000 7.575000 2.250000 ;
        LAYER mcon ;
        RECT 0.675000 1.425000 0.900000 1.650000 ;
        RECT 5.325000 1.950000 5.550000 2.175000 ;
        RECT 6.975000 2.025000 7.200000 2.250000 ;
        LAYER met1 ;
        RECT 0.600000 1.650000 0.975000 1.725000 ;
        RECT 0.600000 1.425000 0.675000 1.650000 ;
        RECT 0.600000 1.350000 0.975000 1.425000 ;
        RECT 0.675000 1.425000 0.900000 1.650000 ;
        RECT 0.900000 1.425000 0.975000 1.650000 ;
        RECT 5.250000 2.175000 5.625000 2.250000 ;
        RECT 5.250000 1.950000 5.325000 2.175000 ;
        RECT 5.250000 1.875000 5.625000 1.950000 ;
        RECT 5.325000 1.950000 5.550000 2.175000 ;
        RECT 6.900000 2.250000 7.275000 2.325000 ;
        RECT 6.900000 2.175000 6.975000 2.250000 ;
        RECT 5.550000 2.025000 6.975000 2.175000 ;
        RECT 5.550000 1.950000 7.275000 2.025000 ;
        RECT 6.975000 2.025000 7.200000 2.250000 ;
        RECT 7.200000 2.025000 7.275000 2.250000 ;
        END
        ANTENNADIFFAREA 2.340000 ;
    END GND
    OBS
        LAYER li ;
        RECT 6.000000 1.350000 8.775000 1.575000 ;
        RECT 1.200000 2.475000 5.775000 2.850000 ;
        RECT 1.200000 2.325000 1.575000 2.475000 ;
        RECT 1.200000 2.100000 1.275000 2.325000 ;
        RECT 1.200000 2.025000 1.575000 2.100000 ;
        RECT 8.775000 1.350000 9.000000 1.575000 ;
        RECT 1.275000 2.100000 1.500000 2.325000 ;
        RECT 6.000000 1.575000 6.300000 1.875000 ;
        RECT 9.000000 1.350000 9.075000 1.575000 ;
        RECT 1.500000 2.100000 1.575000 2.325000 ;
        RECT 8.700000 1.575000 9.075000 1.650000 ;
        RECT 1.800000 3.000000 1.875000 3.225000 ;
        RECT 1.800000 2.850000 2.175000 3.000000 ;
        RECT 1.875000 3.000000 2.100000 3.225000 ;
        RECT 6.000000 1.275000 9.075000 1.350000 ;
        RECT 2.100000 3.000000 2.175000 3.225000 ;
        RECT 6.000000 2.100000 6.300000 3.075000 ;
        RECT 6.000000 1.875000 6.225000 2.100000 ;
        RECT 6.225000 1.875000 6.300000 2.100000 ;
        RECT 7.800000 3.900000 8.025000 4.125000 ;
        RECT 7.800000 3.825000 8.100000 3.900000 ;
        RECT 8.025000 3.900000 8.100000 4.125000 ;
        RECT 5.475000 7.200000 5.850000 7.275000 ;
        RECT 5.475000 6.975000 5.550000 7.200000 ;
        RECT 5.475000 6.900000 5.850000 6.975000 ;
        RECT 5.550000 4.200000 5.775000 6.900000 ;
        RECT 5.550000 4.125000 8.100000 4.200000 ;
        RECT 5.550000 3.975000 7.800000 4.125000 ;
        RECT 5.550000 2.850000 5.775000 3.975000 ;
        RECT 5.550000 6.975000 5.775000 7.200000 ;
        RECT 5.775000 6.975000 5.850000 7.200000 ;
        RECT 6.000000 3.300000 6.300000 3.450000 ;
        RECT 6.000000 3.075000 6.225000 3.300000 ;
        RECT 6.225000 3.075000 6.300000 3.300000 ;
    END
END _0_0std_0_0cells_0_0FAX1

MACRO welltap_svt
    CLASS CORE WELLTAP ;
    FOREIGN welltap_svt 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.200000 BY 2.100000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER li ;
        RECT 0.600000 1.500000 0.900000 1.800000 ;
        END
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER li ;
        RECT 0.600000 0.300000 0.900000 0.600000 ;
        END
    END GND
END welltap_svt

MACRO circuitppnp
   CLASS CORE ;
   FOREIGN circuitppnp 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 432.000000 BY 432.000000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitppnp

MACRO circuitwell
   CLASS CORE ;
   FOREIGN circuitwell 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 432.000000 BY 432.000000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitwell

