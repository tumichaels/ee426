*---------------------------------------------------
* Subcircuit from nor2.ext
*---------------------------------------------------
.subckt nor2 _
* -- connections ---
* -- fets ---
xM1 out in0 a_275_167# Vdd sky130_fd_pr__pfet_01v8  W=0.825 L=0.375
+ AS=0.680625 PS=3.3 AD=0.680625 PD=3.3 nrs=1 nrd=1 nf=1
xM2 GND in0 out Gnd sky130_fd_pr__nfet_01v8 W=0.825 L=0.375
+ AS=0.680625 PS=3.3 AD=1.36125 PD=6.6 nrs=1 nrd=1 nf=1
xM3 a_275_167# in1 Vdd Vdd sky130_fd_pr__pfet_01v8  W=0.825 L=0.375
+ AS=0.680625 PS=3.3 AD=0P PD=0P nrs=1 nrd=1 nf=1
xM4 out in1 GND Gnd sky130_fd_pr__nfet_01v8 W=0.825 L=0.375
+ AS=0P PS=0P AD=0P PD=0P nrs=1 nrd=1 nf=1
* -- caps ---
.ends
*---------------------------------------------------
* Subcircuit from nand2.ext
*---------------------------------------------------
.subckt nand2 _
* -- connections ---
* -- fets ---
xM1 Vdd in0 out Vdd sky130_fd_pr__pfet_01v8  W=0.825 L=0.375
+ AS=0.680625 PS=3.3 AD=1.36125 PD=6.6 nrs=1 nrd=1 nf=1
xM2 out in0 a_85_47# Gnd sky130_fd_pr__nfet_01v8 W=0.825 L=0.375
+ AS=0.680625 PS=3.3 AD=0.680625 PD=3.3 nrs=1 nrd=1 nf=1
xM3 out in1 Vdd Vdd sky130_fd_pr__pfet_01v8  W=0.825 L=0.375
+ AS=0P PS=0P AD=0P PD=0P nrs=1 nrd=1 nf=1
xM4 a_85_47# in1 GND Gnd sky130_fd_pr__nfet_01v8 W=0.825 L=0.375
+ AS=0.680625 PS=3.3 AD=0P PD=0P nrs=1 nrd=1 nf=1
* -- caps ---
.ends
*---------------------------------------------------
* Subcircuit from or4.ext
*---------------------------------------------------
.subckt or4 _
*--- subcircuits ---
xnor2_0 GND nor2
xnor2_1 GND nor2
xnand2_0 GND nand2
* -- connections ---
V1 out xnand2_0:out
V2 in11 xnor2_0:in1
V3 in10 xnor2_0:in0
V4 a_n9_139# xnor2_0:out
V5 xnor2_0:out xnand2_0:in1
V6 a_1_155# xnand2_0:in0
V7 xnand2_0:in0 xnor2_1:out
V8 in00 xnor2_1:in0
V9 in01 xnor2_1:in1
* -- caps ---
.ends
*---------------------------------------------------
* Subcircuit from inv.ext
*---------------------------------------------------
.subckt inv _
* -- connections ---
* -- fets ---
xM1 Vdd in out Vdd sky130_fd_pr__pfet_01v8  W=0.9 L=0.375
+ AS=0.81 PS=3.6 AD=0.81 PD=3.6 nrs=1 nrd=1 nf=1
xM2 GND in out Gnd sky130_fd_pr__nfet_01v8 W=0.9 L=0.375
+ AS=0.81 PS=3.6 AD=0.81 PD=3.6 nrs=1 nrd=1 nf=1
* -- caps ---
.ends
*
*---------------------------------------------------
*  Main extract file or8.ext [scale=1e+06]
*---------------------------------------------------
*
*--- subcircuits ---
xnor2_0 GND nor2
xor4_0 GND or4
xor4_1 GND or4
xinv_0 GND inv
* -- connections ---
V1 in101 xor4_1:in01
V2 m1_30_n6# Vdd
V3 in110 xor4_1:in10
V4 in111 xor4_1:in11
V5 in100 xor4_1:in00
V6 m1_136_n6# Vdd
V7 m1_94_181# GND
V8 GND m1_94_241#
V9 a_42_228# xor4_0:out
V10 xor4_0:out xnor2_0:in0
V11 a_42_212# xor4_1:out
V12 xor4_1:out xnor2_0:in1
V13 m1_30_181# Vdd
V14 Vdd m1_52_209#
V15 a_73_253# xinv_0:in
V16 xinv_0:in xnor2_0:out
V17 in001 xor4_0:in01
V18 in010 xor4_0:in10
V19 out xinv_0:out
V20 in011 xor4_0:in11
V21 in000 xor4_0:in00
* -- caps ---
*--- inferred globals
.global GND
.global Vdd
.global Gnd
