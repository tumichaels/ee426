magic
tech TSMC180
timestamp 1734137093
<< ndiffusion >>
rect 6 21 12 22
rect 6 19 9 21
rect 11 19 12 21
rect 6 12 12 19
rect 14 12 20 22
rect 22 21 28 22
rect 22 19 24 21
rect 26 19 28 21
rect 22 17 28 19
rect 30 20 36 22
rect 30 18 31 20
rect 33 18 36 20
rect 30 17 36 18
rect 22 12 26 17
<< ndcontact >>
rect 9 19 11 21
rect 24 19 26 21
rect 31 18 33 20
<< ntransistor >>
rect 12 12 14 22
rect 20 12 22 22
rect 28 17 30 22
<< pdiffusion >>
rect 6 45 12 46
rect 6 43 9 45
rect 11 43 12 45
rect 6 38 12 43
rect 14 41 20 46
rect 14 39 16 41
rect 18 39 20 41
rect 14 38 20 39
rect 22 45 28 46
rect 22 43 23 45
rect 25 43 28 45
rect 22 38 28 43
rect 30 41 36 46
rect 30 39 31 41
rect 33 39 36 41
rect 30 38 36 39
<< pdcontact >>
rect 9 43 11 45
rect 16 39 18 41
rect 23 43 25 45
rect 31 39 33 41
<< ptransistor >>
rect 12 38 14 46
rect 20 38 22 46
rect 28 38 30 46
<< polysilicon >>
rect 20 57 33 58
rect 6 56 10 57
rect 20 56 30 57
rect 6 54 7 56
rect 9 54 14 56
rect 6 53 14 54
rect 12 46 14 53
rect 20 46 22 56
rect 29 55 30 56
rect 32 55 33 57
rect 29 54 33 55
rect 28 46 30 49
rect 12 22 14 38
rect 20 22 22 38
rect 28 22 30 38
rect 12 9 14 12
rect 20 9 22 12
rect 4 5 8 6
rect 28 5 30 17
rect 4 3 5 5
rect 7 3 30 5
rect 4 2 8 3
<< polycontact >>
rect 7 54 9 56
rect 30 55 32 57
rect 5 3 7 5
<< m1 >>
rect 6 57 9 60
rect 18 57 21 60
rect 30 58 33 60
rect 6 56 10 57
rect 6 54 7 56
rect 9 54 10 56
rect 6 53 10 54
rect 15 54 21 57
rect 29 57 33 58
rect 29 55 30 57
rect 32 55 33 57
rect 29 54 33 55
rect 39 57 45 60
rect 15 50 18 54
rect 9 47 25 50
rect 9 46 12 47
rect 8 45 12 46
rect 8 43 9 45
rect 11 43 12 45
rect 8 42 12 43
rect 22 46 25 47
rect 22 45 26 46
rect 22 43 23 45
rect 25 43 26 45
rect 22 42 26 43
rect 15 41 19 42
rect 15 39 16 41
rect 18 39 19 41
rect 9 36 19 39
rect 30 41 34 42
rect 30 39 31 41
rect 33 39 34 41
rect 30 38 34 39
rect 9 22 12 36
rect 8 21 12 22
rect 8 19 9 21
rect 11 19 12 21
rect 8 18 12 19
rect 22 22 27 23
rect 22 19 23 22
rect 26 19 27 22
rect 22 18 27 19
rect 30 21 33 38
rect 39 23 42 57
rect 37 22 42 23
rect 30 20 34 21
rect 30 18 31 20
rect 33 18 34 20
rect 37 19 38 22
rect 41 19 42 22
rect 37 18 42 19
rect 8 10 11 18
rect 7 9 11 10
rect 5 6 11 9
rect 30 12 34 18
rect 4 5 8 6
rect 4 3 5 5
rect 7 3 8 5
rect 4 2 8 3
rect 30 1 33 12
<< m2c >>
rect 23 21 26 22
rect 23 19 24 21
rect 24 19 26 21
rect 38 19 41 22
<< m2 >>
rect 22 22 42 23
rect 22 19 23 22
rect 26 19 38 22
rect 41 19 42 22
rect 22 18 42 19
<< labels >>
rlabel polysilicon 29 36 29 36 3 _Y
rlabel pdiffusion 31 39 31 39 3 Y
rlabel ndiffusion 23 13 23 13 3 GND
rlabel pdiffusion 23 39 23 39 3 Vdd
rlabel pdiffusion 15 39 15 39 3 _Y
rlabel pdiffusion 7 39 7 39 3 Vdd
rlabel m1 43 58 43 58 3 GND
port 1 e
rlabel m1 7 58 7 58 3 A
port 5 e
rlabel m1 18 57 21 60 5 Vdd
rlabel m1 30 57 33 60 5 B
rlabel m1 31 11 31 11 3 Y
port 4 e
<< end >>
