magic
tech sky130l
timestamp 1731050810
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 28 13 29
rect 8 25 9 28
rect 12 25 13 28
rect 8 19 13 25
rect 15 28 20 29
rect 15 25 16 28
rect 19 25 20 28
rect 15 19 20 25
<< pdc >>
rect 9 25 12 28
rect 16 25 19 28
<< ptransistor >>
rect 13 19 15 29
<< polysilicon >>
rect 13 29 15 31
rect 23 19 28 20
rect 13 17 15 19
rect 23 17 24 19
rect 13 16 24 17
rect 27 16 28 19
rect 13 15 28 16
rect 13 12 15 15
rect 13 4 15 6
<< pc >>
rect 24 16 27 19
<< m1 >>
rect 8 35 12 36
rect 8 32 9 35
rect 9 28 12 32
rect 15 25 16 28
rect 19 25 27 28
rect 9 24 12 25
rect 24 20 27 25
rect 23 19 28 20
rect 23 16 24 19
rect 27 16 28 19
rect 23 15 28 16
rect 9 10 12 11
rect 8 7 9 8
rect 15 8 16 11
rect 19 8 24 11
rect 27 8 28 11
rect 8 4 12 7
rect 23 4 28 8
<< m2c >>
rect 9 32 12 35
rect 24 8 27 11
<< m2 >>
rect 8 35 13 36
rect 8 32 9 35
rect 12 32 13 35
rect 8 31 13 32
rect 23 11 28 12
rect 23 8 24 11
rect 27 8 28 11
rect 23 4 28 8
<< labels >>
rlabel pdiffusion 16 20 16 20 3 x
rlabel polysilicon 14 13 14 13 3 x
rlabel polysilicon 14 18 14 18 3 x
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel m1 9 5 9 5 3 Y
port 2 e
rlabel m1 9 33 9 33 3 Vdd
port 3 e
rlabel m1 21 10 21 10 0 GND
rlabel m2 23 4 28 8 8 GND
<< end >>
