magic
tech sky130l
timestamp 1726527990
<< ndiffusion >>
rect 297 191 308 194
rect 297 186 300 191
rect 305 186 308 191
rect 297 183 308 186
rect 297 175 308 178
rect 297 170 300 175
rect 305 170 308 175
rect 297 167 308 170
rect 297 159 308 162
rect 297 154 300 159
rect 305 154 308 159
rect 297 151 308 154
<< ndc >>
rect 300 186 305 191
rect 300 170 305 175
rect 300 154 305 159
<< ntransistor >>
rect 297 178 308 183
rect 297 162 308 167
<< pdiffusion >>
rect 275 191 286 194
rect 275 186 278 191
rect 283 186 286 191
rect 275 183 286 186
rect 275 167 286 178
rect 275 159 286 162
rect 275 154 278 159
rect 283 154 286 159
rect 275 151 286 154
<< pdc >>
rect 278 186 283 191
rect 278 154 283 159
<< ptransistor >>
rect 275 178 286 183
rect 275 162 286 167
<< polysilicon >>
rect 256 178 275 183
rect 286 178 297 183
rect 308 178 310 183
rect 256 162 275 167
rect 286 162 297 167
rect 308 162 310 167
<< m1 >>
rect 288 192 295 194
rect 277 191 295 192
rect 277 186 278 191
rect 283 186 295 191
rect 277 185 295 186
rect 299 191 316 192
rect 299 186 300 191
rect 305 186 316 191
rect 299 185 316 186
rect 288 176 295 185
rect 288 175 306 176
rect 288 170 300 175
rect 305 170 306 175
rect 288 169 306 170
rect 309 160 316 185
rect 267 159 284 160
rect 267 154 278 159
rect 283 154 284 159
rect 267 153 284 154
rect 299 159 316 160
rect 299 154 300 159
rect 305 154 316 159
rect 299 153 316 154
<< labels >>
rlabel m1 309 153 316 192 3 GND!
rlabel m1 288 169 295 194 1 out
rlabel polysilicon 256 178 275 183 7 in0
rlabel polysilicon 256 162 275 167 7 in1
rlabel m1 267 153 278 160 7 Vdd!
<< end >>
