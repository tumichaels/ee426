*
*---------------------------------------------------
*  Main extract file inv.ext [scale=1e+06]
*---------------------------------------------------
*
* -- connections ---
* -- fets ---
xM1 Vdd in out Vdd sky130_fd_pr__pfet_01v8  W=0.9 L=0.375
+ AS=0.81 PS=3.6 AD=0.81 PD=3.6 nrs=1 nrd=1 nf=1
xM2 GND in out Gnd sky130_fd_pr__nfet_01v8 W=0.9 L=0.375
+ AS=0.81 PS=3.6 AD=0.81 PD=3.6 nrs=1 nrd=1 nf=1
* -- caps ---
*--- inferred globals
.global Vdd
.global GND
.global Gnd
