magic
tech sky130l
timestamp 1731041397
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
rect 22 10 27 12
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 12
rect 20 6 22 12
<< pdiffusion >>
rect 8 33 13 34
rect 8 30 9 33
rect 12 30 13 33
rect 8 19 13 30
rect 15 19 20 34
rect 22 23 27 34
rect 22 20 23 23
rect 26 20 27 23
rect 22 19 27 20
<< pdc >>
rect 9 30 12 33
rect 23 20 26 23
<< ptransistor >>
rect 13 19 15 34
rect 20 19 22 34
<< polysilicon >>
rect 15 44 20 45
rect 15 42 16 44
rect 13 41 16 42
rect 19 41 20 44
rect 13 40 20 41
rect 13 34 15 40
rect 20 34 22 36
rect 30 34 35 35
rect 30 31 31 34
rect 34 31 35 34
rect 30 30 35 31
rect 13 12 15 19
rect 20 17 22 19
rect 32 17 34 30
rect 20 15 34 17
rect 20 12 22 15
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 16 41 19 44
rect 31 31 34 34
<< m1 >>
rect 16 44 20 45
rect 8 39 12 44
rect 8 36 9 39
rect 19 41 20 44
rect 16 36 20 41
rect 32 39 36 45
rect 31 36 36 39
rect 9 33 12 36
rect 31 34 34 36
rect 31 30 34 31
rect 9 29 12 30
rect 23 23 26 24
rect 23 16 26 20
rect 9 13 26 16
rect 9 10 12 13
rect 23 10 26 13
rect 8 7 9 8
rect 15 7 16 10
rect 19 7 20 10
rect 8 4 12 7
rect 23 6 26 7
rect 35 5 36 8
rect 32 4 36 5
<< m2c >>
rect 9 36 12 39
rect 16 7 19 10
rect 32 5 35 8
<< m2 >>
rect 8 40 12 44
rect 8 39 13 40
rect 8 36 9 39
rect 12 36 13 39
rect 8 35 13 36
rect 15 10 20 11
rect 15 7 16 10
rect 19 9 34 10
rect 19 8 36 9
rect 19 7 20 8
rect 15 6 20 7
rect 31 5 32 8
rect 35 5 36 8
rect 31 4 36 5
<< labels >>
rlabel space 0 0 40 48 6 prboundary
rlabel polysilicon 35 32 35 32 3 B
rlabel polysilicon 33 18 33 18 3 B
rlabel ndiffusion 27 8 27 8 3 Y
rlabel polysilicon 31 31 31 31 3 B
rlabel polysilicon 31 32 31 32 3 B
rlabel polysilicon 31 35 31 35 3 B
rlabel pdiffusion 27 21 27 21 3 Y
rlabel ndiffusion 23 7 23 7 3 Y
rlabel ndiffusion 23 8 23 8 3 Y
rlabel ndiffusion 23 11 23 11 3 Y
rlabel pdiffusion 23 20 23 20 3 Y
rlabel pdiffusion 23 21 23 21 3 Y
rlabel pdiffusion 23 24 23 24 3 Y
rlabel polysilicon 21 5 21 5 3 B
rlabel ntransistor 21 7 21 7 3 B
rlabel polysilicon 21 13 21 13 3 B
rlabel polysilicon 21 16 21 16 3 B
rlabel polysilicon 21 18 21 18 3 B
rlabel ptransistor 21 20 21 20 3 B
rlabel polysilicon 21 35 21 35 3 B
rlabel ndiffusion 13 8 13 8 3 Y
rlabel pdiffusion 13 31 13 31 3 Vdd
rlabel polysilicon 16 43 16 43 3 A
rlabel polysilicon 16 45 16 45 3 A
rlabel polysilicon 14 5 14 5 3 A
rlabel ntransistor 14 7 14 7 3 A
rlabel polysilicon 14 13 14 13 3 A
rlabel ptransistor 14 20 14 20 3 A
rlabel polysilicon 14 35 14 35 3 A
rlabel polysilicon 14 41 14 41 3 A
rlabel polysilicon 14 42 14 42 3 A
rlabel ndiffusion 9 7 9 7 3 Y
rlabel ndiffusion 9 11 9 11 3 Y
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel pdiffusion 9 31 9 31 3 Vdd
rlabel pdiffusion 9 34 9 34 3 Vdd
rlabel m1 33 40 33 40 3 B
port 1 e
rlabel m1 32 31 32 31 3 B
port 1 e
rlabel pc 32 32 32 32 3 B
port 1 e
rlabel m1 32 35 32 35 3 B
port 1 e
rlabel m1 32 37 32 37 3 B
port 1 e
rlabel ndc 24 8 24 8 3 Y
port 2 e
rlabel m1 24 11 24 11 3 Y
port 2 e
rlabel m1 24 17 24 17 3 Y
port 2 e
rlabel pdc 24 21 24 21 3 Y
port 2 e
rlabel m1 24 24 24 24 3 Y
port 2 e
rlabel m1 20 42 20 42 3 A
port 3 e
rlabel m1 33 5 33 5 3 GND
rlabel m1 17 37 17 37 3 A
port 3 e
rlabel pc 17 42 17 42 3 A
port 3 e
rlabel m1 17 45 17 45 3 A
port 3 e
rlabel m1 24 7 24 7 3 Y
port 2 e
rlabel ndc 10 8 10 8 3 Y
port 2 e
rlabel m1 10 11 10 11 3 Y
port 2 e
rlabel m1 10 14 10 14 3 Y
port 2 e
rlabel m1 10 30 10 30 3 Vdd
rlabel pdc 10 31 10 31 3 Vdd
rlabel m1 10 34 10 34 3 Vdd
rlabel m1 9 5 9 5 3 Y
port 2 e
rlabel m1 9 8 9 8 3 Y
port 2 e
rlabel m2 36 6 36 6 3 GND
rlabel m2c 33 6 33 6 3 GND
rlabel m2 32 5 32 5 3 GND
rlabel m2 32 6 32 6 3 GND
rlabel m2 20 8 20 8 3 GND
rlabel m2 20 9 20 9 3 GND
rlabel m2 20 10 20 10 3 GND
rlabel m2c 17 8 17 8 3 GND
rlabel m2 16 7 16 7 3 GND
rlabel m2 16 8 16 8 3 GND
rlabel m2 16 11 16 11 3 GND
rlabel m2 13 37 13 37 3 Vdd
rlabel m2c 10 37 10 37 3 Vdd
rlabel m2 9 36 9 36 3 Vdd
rlabel m2 9 37 9 37 3 Vdd
rlabel m2 9 40 9 40 3 Vdd
rlabel m2 9 41 9 41 3 Vdd
<< end >>
