magic
tech sky130l
timestamp 1730908935
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 10 20 12
rect 15 7 16 10
rect 19 7 20 10
rect 15 6 20 7
<< ndc >>
rect 9 7 12 10
rect 16 7 19 10
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 23 13 27
rect 8 20 9 23
rect 12 20 13 23
rect 8 19 13 20
rect 15 23 20 27
rect 15 20 16 23
rect 19 20 20 23
rect 15 19 20 20
<< pdc >>
rect 9 20 12 23
rect 16 20 19 23
<< ptransistor >>
rect 13 19 15 27
<< polysilicon >>
rect 13 27 15 29
rect 13 17 15 19
rect 23 17 28 18
rect 13 15 24 17
rect 13 12 15 15
rect 23 14 24 15
rect 27 14 28 17
rect 23 13 28 14
rect 13 4 15 6
<< pc >>
rect 24 14 27 17
<< m1 >>
rect 8 31 12 32
rect 8 28 9 31
rect 16 28 20 32
rect 24 28 28 32
rect 9 23 12 24
rect 16 23 19 28
rect 15 20 16 23
rect 19 20 20 23
rect 9 10 12 20
rect 23 17 28 18
rect 19 14 24 17
rect 27 14 28 17
rect 23 13 28 14
rect 8 7 9 8
rect 8 4 12 7
rect 16 10 19 11
rect 16 6 19 7
<< m2c >>
rect 9 28 12 31
rect 24 25 27 28
rect 16 14 19 17
rect 16 7 19 10
<< m2 >>
rect 8 31 13 32
rect 8 28 9 31
rect 12 28 13 31
rect 8 27 13 28
rect 11 17 13 27
rect 23 28 28 29
rect 23 25 24 28
rect 27 25 28 28
rect 23 24 28 25
rect 15 17 20 18
rect 11 15 16 17
rect 15 14 16 15
rect 19 14 20 17
rect 15 13 20 14
rect 15 10 20 11
rect 23 10 25 24
rect 15 7 16 10
rect 19 8 25 10
rect 19 7 20 8
rect 15 6 20 7
<< labels >>
rlabel space 0 0 32 36 6 prboundary
rlabel polysilicon 24 15 24 15 3 A
rlabel ndiffusion 13 8 13 8 3 Y
rlabel pdiffusion 16 20 16 20 3 Vdd
rlabel pdiffusion 16 24 16 24 3 Vdd
rlabel pdiffusion 13 21 13 21 3 Y
rlabel polysilicon 14 5 14 5 3 A
rlabel ntransistor 14 7 14 7 3 A
rlabel polysilicon 14 13 14 13 3 A
rlabel polysilicon 14 16 14 16 3 A
rlabel polysilicon 14 18 14 18 3 A
rlabel ptransistor 14 20 14 20 3 A
rlabel polysilicon 14 28 14 28 3 A
rlabel ndiffusion 9 7 9 7 3 Y
rlabel ndiffusion 9 11 9 11 3 Y
rlabel pdiffusion 9 20 9 20 3 Y
rlabel pdiffusion 9 21 9 21 3 Y
rlabel pdiffusion 9 24 9 24 3 Y
rlabel m1 28 15 28 15 3 A
port 1 e
rlabel m1 24 14 24 14 3 A
port 1 e
rlabel pc 25 15 25 15 3 A
port 1 e
rlabel m1 24 18 24 18 3 A
port 1 e
rlabel m1 25 29 25 29 3 GND
rlabel m1 20 21 20 21 3 Vdd
rlabel m1 17 11 17 11 3 GND
rlabel pdc 17 21 17 21 3 Vdd
rlabel m1 17 24 17 24 3 Vdd
rlabel m1 17 29 17 29 3 Vdd
rlabel m1 16 21 16 21 3 Vdd
rlabel m1 17 7 17 7 3 GND
rlabel ndc 10 8 10 8 3 Y
port 2 e
rlabel m1 10 11 10 11 3 Y
port 2 e
rlabel pdc 10 21 10 21 3 Y
port 2 e
rlabel m1 10 24 10 24 3 Y
port 2 e
rlabel m1 9 5 9 5 3 Y
port 2 e
rlabel m1 9 8 9 8 3 Y
port 2 e
rlabel m2 28 26 28 26 3 GND
rlabel m2c 25 26 25 26 3 GND
rlabel m2 24 25 24 25 3 GND
rlabel m2 24 26 24 26 3 GND
rlabel m2 20 8 20 8 3 GND
rlabel m2 20 9 20 9 3 GND
rlabel m2 24 11 24 11 3 GND
rlabel m2 20 15 20 15 3 A
port 1 e
rlabel m2c 17 8 17 8 3 GND
rlabel m2c 17 15 17 15 3 A
port 1 e
rlabel m2 16 18 16 18 3 A
port 1 e
rlabel m2 24 29 24 29 3 GND
rlabel m2 16 7 16 7 3 GND
rlabel m2 16 8 16 8 3 GND
rlabel m2 16 11 16 11 3 GND
rlabel m2 16 14 16 14 3 A
port 1 e
rlabel m2 16 15 16 15 3 A
port 1 e
rlabel m2 12 16 12 16 3 A
port 1 e
rlabel m2 12 18 12 18 3 A
port 1 e
rlabel m2 13 29 13 29 3 A
port 1 e
rlabel m2c 10 29 10 29 3 A
port 1 e
rlabel m2 9 28 9 28 3 A
port 1 e
rlabel m2 9 29 9 29 3 A
port 1 e
rlabel m2 9 32 9 32 3 A
port 1 e
<< end >>
