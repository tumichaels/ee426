magic
tech TSMC180
timestamp 1734150867
<< ndiffusion >>
rect 6 10 12 12
rect 6 8 8 10
rect 10 8 12 10
rect 6 7 12 8
rect 14 7 20 12
rect 22 10 28 12
rect 22 8 24 10
rect 26 8 28 10
rect 22 7 28 8
<< ndcontact >>
rect 8 8 10 10
rect 24 8 26 10
<< ntransistor >>
rect 12 7 14 12
rect 20 7 22 12
<< pdiffusion >>
rect 6 42 12 43
rect 6 40 7 42
rect 9 40 12 42
rect 6 28 12 40
rect 14 28 20 43
rect 22 32 28 43
rect 22 30 25 32
rect 27 30 28 32
rect 22 28 28 30
<< pdcontact >>
rect 7 40 9 42
rect 25 30 27 32
<< ptransistor >>
rect 12 28 14 43
rect 20 28 22 43
<< polysilicon >>
rect 18 57 22 58
rect 18 55 19 57
rect 21 55 22 57
rect 18 54 22 55
rect 12 49 16 50
rect 12 47 13 49
rect 15 47 16 49
rect 12 46 16 47
rect 12 43 14 46
rect 20 43 22 54
rect 12 12 14 28
rect 20 12 22 28
rect 12 4 14 7
rect 20 4 22 7
<< polycontact >>
rect 19 55 21 57
rect 13 47 15 49
<< m1 >>
rect 6 43 9 64
rect 12 50 15 64
rect 18 58 21 64
rect 18 57 22 58
rect 18 55 19 57
rect 21 55 22 57
rect 18 54 22 55
rect 12 49 16 50
rect 12 47 13 49
rect 15 47 16 49
rect 12 46 16 47
rect 25 43 28 64
rect 6 42 10 43
rect 6 40 7 42
rect 9 40 10 42
rect 6 39 10 40
rect 24 32 28 43
rect 24 30 25 32
rect 27 30 28 32
rect 24 28 28 30
rect 15 24 28 28
rect 7 10 11 11
rect 7 8 8 10
rect 10 8 11 10
rect 15 9 19 24
rect 23 10 27 11
rect 7 6 11 8
rect 23 8 24 10
rect 26 8 27 10
rect 23 6 27 8
rect 7 3 27 6
rect 24 -4 27 3
<< labels >>
rlabel pdiffusion 23 29 23 29 3 Y
rlabel polysilicon 21 13 21 13 3 B
rlabel polysilicon 21 26 21 26 3 B
rlabel ndiffusion 15 8 15 8 3 Y
rlabel polysilicon 13 13 13 13 3 A
rlabel polysilicon 13 26 13 26 3 A
rlabel pdiffusion 7 29 7 29 3 Vdd
rlabel m1 19 55 19 55 3 B
port 3 e
rlabel m1 13 55 13 55 3 A
port 5 e
rlabel m1 7 55 7 55 3 Vdd
port 2 e
rlabel m1 26 2 26 2 3 GND
port 1 e
rlabel m1 26 55 26 55 3 Y
port 4 e
rlabel ndiffusion 7 8 7 8 3 GND
rlabel ndiffusion 23 8 23 8 3 GND
<< end >>
