magic
tech sky130l
timestamp 1731048377
<< ndiffusion >>
rect 8 10 13 16
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 15 20 16
rect 15 12 16 15
rect 19 12 20 15
rect 15 6 20 12
rect 22 10 27 16
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
<< ndc >>
rect 9 7 12 10
rect 16 12 19 15
rect 23 7 26 10
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
<< pdiffusion >>
rect 8 48 13 53
rect 8 43 9 48
rect 12 43 13 48
rect 8 23 13 43
rect 15 23 20 53
rect 22 32 27 53
rect 22 26 23 32
rect 26 26 27 32
rect 22 23 27 26
<< pdc >>
rect 9 43 12 48
rect 23 26 26 32
<< ptransistor >>
rect 13 23 15 53
rect 20 23 22 53
<< polysilicon >>
rect 8 61 15 62
rect 8 58 9 61
rect 12 58 15 61
rect 8 57 15 58
rect 13 53 15 57
rect 20 61 28 62
rect 20 58 24 61
rect 27 58 28 61
rect 20 57 28 58
rect 20 53 22 57
rect 13 16 15 23
rect 20 16 22 23
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 9 58 12 61
rect 24 58 27 61
<< m1 >>
rect 8 62 12 68
rect 16 67 20 68
rect 16 64 17 67
rect 8 61 13 62
rect 8 58 9 61
rect 12 58 13 61
rect 8 57 13 58
rect 8 48 13 49
rect 8 43 9 48
rect 12 46 13 48
rect 16 46 20 64
rect 24 62 28 68
rect 23 61 28 62
rect 23 58 24 61
rect 27 58 28 61
rect 23 57 28 58
rect 12 43 20 46
rect 8 42 20 43
rect 22 32 27 33
rect 22 26 23 32
rect 26 26 27 32
rect 22 22 27 26
rect 15 21 27 22
rect 15 17 36 21
rect 15 15 20 17
rect 15 12 16 15
rect 19 12 20 15
rect 9 10 12 11
rect 8 7 9 8
rect 23 10 27 11
rect 22 8 23 9
rect 12 7 23 8
rect 26 7 27 10
rect 8 6 26 7
rect 8 5 25 6
rect 8 4 13 5
rect 32 4 36 17
<< m2c >>
rect 17 64 20 67
rect 9 7 12 10
<< m2 >>
rect 16 67 21 68
rect 16 64 17 67
rect 20 64 21 67
rect 16 63 21 64
rect 8 10 13 11
rect 8 7 9 10
rect 12 7 13 10
rect 8 4 13 7
<< labels >>
rlabel m1 9 65 9 65 3 A
port 5 e
rlabel m1 25 65 25 65 3 B
port 2 e
rlabel m1 17 65 17 65 3 Vdd
port 3 e
rlabel m1 33 5 33 5 3 Y
port 1 e
rlabel m2 8 4 13 7 2 GND
<< end >>
