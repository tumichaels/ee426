magic
tech sky130l
timestamp 1730909060
<< ndiffusion >>
rect 8 10 13 12
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 11 20 12
rect 15 8 16 11
rect 19 8 20 11
rect 15 6 20 8
<< ndc >>
rect 9 7 12 10
rect 16 8 19 11
<< ntransistor >>
rect 13 6 15 12
<< pdiffusion >>
rect 8 28 13 29
rect 8 25 9 28
rect 12 25 13 28
rect 8 19 13 25
rect 15 28 20 29
rect 15 25 16 28
rect 19 25 20 28
rect 15 19 20 25
<< pdc >>
rect 9 25 12 28
rect 16 25 19 28
<< ptransistor >>
rect 13 19 15 29
<< polysilicon >>
rect 13 29 15 31
rect 23 19 28 20
rect 13 17 15 19
rect 23 17 24 19
rect 13 16 24 17
rect 27 16 28 19
rect 13 15 28 16
rect 13 12 15 15
rect 13 4 15 6
<< pc >>
rect 24 16 27 19
<< m1 >>
rect 8 32 12 36
rect 9 28 12 32
rect 23 35 28 36
rect 23 32 24 35
rect 27 32 28 35
rect 23 31 28 32
rect 15 25 16 28
rect 19 25 27 28
rect 9 24 12 25
rect 24 20 27 25
rect 23 19 28 20
rect 23 16 24 19
rect 27 16 28 19
rect 23 15 28 16
rect 9 10 12 11
rect 8 7 9 8
rect 15 8 16 11
rect 19 8 24 11
rect 8 4 12 7
<< m2c >>
rect 24 32 27 35
rect 24 8 27 11
<< m2 >>
rect 23 35 28 36
rect 23 32 24 35
rect 27 32 28 35
rect 23 31 28 32
rect 24 12 27 31
rect 23 11 28 12
rect 23 8 24 11
rect 27 8 28 11
rect 23 7 28 8
<< labels >>
rlabel space 0 0 32 40 6 prboundary
rlabel polysilicon 24 18 24 18 3 x
rlabel ndiffusion 16 7 16 7 3 GND
rlabel ndiffusion 16 12 16 12 3 GND
rlabel ndiffusion 13 8 13 8 3 Y
rlabel pdiffusion 16 20 16 20 3 x
rlabel pdiffusion 16 29 16 29 3 x
rlabel pdiffusion 13 26 13 26 3 Vdd
rlabel polysilicon 14 5 14 5 3 x
rlabel ntransistor 14 7 14 7 3 x
rlabel polysilicon 14 13 14 13 3 x
rlabel polysilicon 14 16 14 16 3 x
rlabel polysilicon 14 17 14 17 3 x
rlabel polysilicon 14 18 14 18 3 x
rlabel ptransistor 14 20 14 20 3 x
rlabel polysilicon 14 30 14 30 3 x
rlabel ndiffusion 9 7 9 7 3 Y
rlabel ndiffusion 9 11 9 11 3 Y
rlabel pdiffusion 9 20 9 20 3 Vdd
rlabel pdiffusion 9 26 9 26 3 Vdd
rlabel pdiffusion 9 29 9 29 3 Vdd
rlabel m1 28 17 28 17 3 x
rlabel pc 25 17 25 17 3 x
rlabel m1 25 21 25 21 3 x
rlabel m1 24 16 24 16 3 x
rlabel m1 24 17 24 17 3 x
rlabel m1 24 20 24 20 3 x
rlabel m1 20 9 20 9 3 GND
rlabel m1 20 26 20 26 3 x
rlabel ndc 17 9 17 9 3 GND
rlabel pdc 17 26 17 26 3 x
rlabel m1 16 9 16 9 3 GND
rlabel m1 16 26 16 26 3 x
rlabel ndc 10 8 10 8 3 Y
port 1 e
rlabel m1 10 11 10 11 3 Y
port 1 e
rlabel m1 10 25 10 25 3 Vdd
rlabel pdc 10 26 10 26 3 Vdd
rlabel m1 10 29 10 29 3 Vdd
rlabel m1 9 5 9 5 3 Y
port 1 e
rlabel m1 9 8 9 8 3 Y
port 1 e
rlabel m1 9 33 9 33 3 Vdd
rlabel m2 28 9 28 9 3 GND
rlabel m2 28 33 28 33 3 GND
rlabel m2c 25 9 25 9 3 GND
rlabel m2 25 13 25 13 3 GND
rlabel m2c 25 33 25 33 3 GND
rlabel m2 24 8 24 8 3 GND
rlabel m2 24 9 24 9 3 GND
rlabel m2 24 12 24 12 3 GND
rlabel m2 24 32 24 32 3 GND
rlabel m2 24 33 24 33 3 GND
rlabel m2 24 36 24 36 3 GND
<< end >>
