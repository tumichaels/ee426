magic
tech TSMC180
timestamp 1734135876
<< ndiffusion >>
rect 6 21 12 22
rect 6 19 7 21
rect 9 19 12 21
rect 25 19 29 22
rect 31 19 39 22
rect 6 18 10 19
rect 35 13 39 19
rect 35 11 36 13
rect 38 11 39 13
rect 35 7 39 11
rect 41 7 45 22
rect 47 7 51 22
rect 53 21 59 22
rect 53 19 54 21
rect 56 19 59 21
rect 53 16 59 19
rect 63 21 69 22
rect 63 19 64 21
rect 66 19 69 21
rect 63 16 69 19
rect 53 7 57 16
<< ndcontact >>
rect 7 19 9 21
rect 36 11 38 13
rect 54 19 56 21
rect 64 19 66 21
<< ntransistor >>
rect 12 19 25 22
rect 29 19 31 22
rect 39 7 41 22
rect 45 7 47 22
rect 51 7 53 22
rect 59 16 63 22
<< pdiffusion >>
rect 6 41 10 42
rect 35 41 39 56
rect 6 39 7 41
rect 9 39 12 41
rect 6 38 12 39
rect 18 38 29 41
rect 31 39 36 41
rect 38 39 39 41
rect 31 38 39 39
rect 41 38 45 56
rect 47 38 51 56
rect 53 54 57 56
rect 53 52 54 54
rect 56 52 57 54
rect 53 44 57 52
rect 53 38 59 44
rect 63 41 69 44
rect 63 39 64 41
rect 66 39 69 41
rect 63 38 69 39
<< pdcontact >>
rect 7 39 9 41
rect 36 39 38 41
rect 54 52 56 54
rect 64 39 66 41
<< ptransistor >>
rect 12 38 18 41
rect 29 38 31 41
rect 39 38 41 56
rect 45 38 47 56
rect 51 38 53 56
rect 59 38 63 44
<< polysilicon >>
rect 18 67 22 68
rect 18 65 19 67
rect 21 66 22 67
rect 21 65 47 66
rect 18 64 47 65
rect 6 62 10 63
rect 6 60 7 62
rect 9 60 10 62
rect 6 59 41 60
rect 7 58 41 59
rect 39 56 41 58
rect 45 56 47 64
rect 51 63 55 64
rect 51 61 52 63
rect 54 61 55 63
rect 51 60 55 61
rect 51 56 53 60
rect 13 47 18 48
rect 13 44 14 47
rect 17 44 18 47
rect 28 47 32 48
rect 28 45 29 47
rect 31 45 32 47
rect 28 44 32 45
rect 12 41 18 44
rect 29 41 31 44
rect 59 44 63 47
rect 12 35 18 38
rect 13 28 18 29
rect 13 25 14 28
rect 17 25 18 28
rect 12 22 25 25
rect 29 22 31 38
rect 39 22 41 38
rect 45 22 47 38
rect 51 22 53 38
rect 59 22 63 38
rect 12 16 25 19
rect 29 16 31 19
rect 59 14 63 16
rect 59 13 64 14
rect 59 10 60 13
rect 63 10 64 13
rect 59 9 64 10
rect 39 4 41 7
rect 45 4 47 7
rect 51 4 53 7
<< polycontact >>
rect 19 65 21 67
rect 7 60 9 62
rect 52 61 54 63
rect 14 44 17 47
rect 29 45 31 47
rect 14 25 17 28
rect 60 10 63 13
<< m1 >>
rect 6 63 9 76
rect 18 68 21 76
rect 18 67 22 68
rect 18 65 19 67
rect 21 65 22 67
rect 18 64 22 65
rect 36 64 39 76
rect 36 63 55 64
rect 6 62 10 63
rect 6 60 7 62
rect 9 60 10 62
rect 36 61 52 63
rect 54 61 55 63
rect 51 60 55 61
rect 6 59 10 60
rect 52 55 57 56
rect 60 55 63 76
rect 52 54 63 55
rect 7 52 54 54
rect 56 52 63 54
rect 7 51 63 52
rect 7 42 10 51
rect 13 47 18 48
rect 13 44 14 47
rect 17 46 18 47
rect 28 47 67 48
rect 17 44 24 46
rect 28 45 29 47
rect 31 45 67 47
rect 28 44 32 45
rect 13 43 24 44
rect 6 41 10 42
rect 6 39 7 41
rect 9 39 10 41
rect 6 38 10 39
rect 7 29 10 38
rect 7 28 18 29
rect 7 26 14 28
rect 13 25 14 26
rect 17 25 18 28
rect 13 24 18 25
rect 6 21 10 22
rect 21 21 24 43
rect 64 42 67 45
rect 35 41 39 42
rect 35 39 36 41
rect 38 39 39 41
rect 35 38 39 39
rect 28 21 33 22
rect 6 19 7 21
rect 9 19 29 21
rect 6 18 29 19
rect 32 18 33 21
rect 28 17 33 18
rect 36 14 39 38
rect 63 41 67 42
rect 63 39 64 41
rect 66 39 67 41
rect 63 38 67 39
rect 63 22 66 38
rect 72 22 75 28
rect 52 21 57 22
rect 52 18 53 21
rect 56 18 57 21
rect 63 21 67 22
rect 63 19 64 21
rect 66 19 67 21
rect 63 18 67 19
rect 70 21 75 22
rect 70 18 71 21
rect 74 18 75 21
rect 52 17 57 18
rect 70 17 75 18
rect 35 13 64 14
rect 3 11 36 13
rect 38 11 60 13
rect 3 10 39 11
rect 59 10 60 11
rect 63 10 64 13
rect 3 7 9 10
rect 59 9 64 10
rect 6 3 9 7
rect 5 -1 10 3
<< m2c >>
rect 29 18 32 21
rect 53 19 54 21
rect 54 19 56 21
rect 53 18 56 19
rect 71 18 74 21
<< m2 >>
rect 28 21 75 22
rect 28 18 29 21
rect 32 18 53 21
rect 56 18 71 21
rect 74 18 75 21
rect 28 17 75 18
<< labels >>
rlabel ndiffusion 54 8 54 8 3 GND
rlabel polysilicon 30 23 30 23 3 #10
rlabel polysilicon 30 36 30 36 3 #10
rlabel polysilicon 13 23 13 23 3 Vdd
rlabel polysilicon 13 36 13 36 3 GND
rlabel m1 61 68 61 68 3 Vdd
port 8 e
rlabel m1 18 67 21 70 5 in(1)
rlabel m1 7 11 7 11 3 out
port 11 e
rlabel m1 7 68 7 68 3 in(0)
port 12 e
rlabel m1 37 68 37 68 3 in(2)
port 9 e
rlabel m1 6 7 9 13 3 out
rlabel m1 72 22 75 28 7 GND
<< end >>
