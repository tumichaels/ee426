magic
tech sky130l
timestamp 1726527220
<< ndiffusion >>
rect 85 71 96 74
rect 85 66 88 71
rect 93 66 96 71
rect 85 63 96 66
rect 85 47 96 58
rect 85 39 96 42
rect 85 34 88 39
rect 93 34 96 39
rect 85 31 96 34
<< ndc >>
rect 88 66 93 71
rect 88 34 93 39
<< ntransistor >>
rect 85 58 96 63
rect 85 42 96 47
<< pdiffusion >>
rect 63 71 74 74
rect 63 66 66 71
rect 71 66 74 71
rect 63 63 74 66
rect 63 55 74 58
rect 63 50 66 55
rect 71 50 74 55
rect 63 47 74 50
rect 63 39 74 42
rect 63 34 66 39
rect 71 34 74 39
rect 63 31 74 34
<< pdc >>
rect 66 66 71 71
rect 66 50 71 55
rect 66 34 71 39
<< ptransistor >>
rect 63 58 74 63
rect 63 42 74 47
<< polysilicon >>
rect 44 58 63 63
rect 74 58 85 63
rect 96 58 98 63
rect 44 42 63 47
rect 74 42 85 47
rect 96 42 98 47
<< m1 >>
rect 76 72 83 74
rect 55 71 72 72
rect 55 66 66 71
rect 71 66 72 71
rect 55 65 72 66
rect 76 71 94 72
rect 76 66 88 71
rect 93 66 94 71
rect 76 65 94 66
rect 55 40 62 65
rect 76 56 83 65
rect 65 55 83 56
rect 65 50 66 55
rect 71 50 83 55
rect 65 49 83 50
rect 55 39 72 40
rect 55 34 66 39
rect 71 34 72 39
rect 55 33 72 34
rect 87 39 104 40
rect 87 34 88 39
rect 93 34 104 39
rect 87 33 104 34
<< labels >>
rlabel m1 55 33 62 72 7 Vdd!
rlabel m1 76 49 83 74 1 out
rlabel m1 93 33 104 40 3 GND!
rlabel polysilicon 44 58 63 63 7 in0
rlabel polysilicon 44 42 63 47 7 in1
<< end >>
