magic
tech sky130l
timestamp 1731009272
<< ndiffusion >>
rect 8 12 13 16
rect 8 8 9 12
rect 12 8 13 12
rect 8 6 13 8
rect 15 15 20 16
rect 15 12 16 15
rect 19 12 20 15
rect 15 6 20 12
rect 22 12 27 16
rect 22 8 23 12
rect 26 8 27 12
rect 22 6 27 8
<< ndc >>
rect 9 8 12 12
rect 16 12 19 15
rect 23 8 26 12
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
<< pdiffusion >>
rect 8 48 13 53
rect 8 43 9 48
rect 12 43 13 48
rect 8 23 13 43
rect 15 23 20 53
rect 22 32 27 53
rect 22 26 23 32
rect 26 26 27 32
rect 22 23 27 26
<< pdc >>
rect 9 43 12 48
rect 23 26 26 32
<< ptransistor >>
rect 13 23 15 53
rect 20 23 22 53
<< polysilicon >>
rect 8 61 15 62
rect 8 58 9 61
rect 12 58 15 61
rect 8 57 15 58
rect 13 53 15 57
rect 20 61 28 62
rect 20 58 24 61
rect 27 58 28 61
rect 20 57 28 58
rect 20 53 22 57
rect 13 16 15 23
rect 20 16 22 23
rect 13 4 15 6
rect 20 4 22 6
<< pc >>
rect 9 58 12 61
rect 24 58 27 61
<< m1 >>
rect 8 62 12 68
rect 8 61 13 62
rect 8 58 9 61
rect 12 58 13 61
rect 8 57 13 58
rect 8 48 13 49
rect 8 43 9 48
rect 12 46 13 48
rect 16 46 20 68
rect 24 62 28 68
rect 23 61 28 62
rect 23 58 24 61
rect 27 58 28 61
rect 23 57 28 58
rect 12 43 20 46
rect 8 42 20 43
rect 22 32 27 33
rect 22 26 23 32
rect 26 26 27 32
rect 22 22 27 26
rect 15 21 27 22
rect 32 21 36 68
rect 15 17 36 21
rect 15 15 20 17
rect 8 12 12 13
rect 8 8 9 12
rect 15 12 16 15
rect 19 12 20 15
rect 15 11 20 12
rect 23 12 27 13
rect 26 8 27 12
rect 8 4 27 8
<< labels >>
rlabel space 0 0 40 72 6 prboundary
rlabel ndiffusion 23 7 23 7 3 GND
rlabel ndiffusion 23 9 23 9 3 GND
rlabel ndiffusion 23 13 23 13 3 GND
rlabel pdiffusion 23 24 23 24 3 Y
rlabel polysilicon 21 5 21 5 3 B
rlabel ntransistor 21 7 21 7 3 B
rlabel polysilicon 21 17 21 17 3 B
rlabel ptransistor 21 24 21 24 3 B
rlabel polysilicon 21 54 21 54 3 B
rlabel polysilicon 21 58 21 58 3 B
rlabel polysilicon 21 59 21 59 3 B
rlabel polysilicon 21 62 21 62 3 B
rlabel ndiffusion 16 7 16 7 3 Y
rlabel ndiffusion 13 9 13 9 3 GND
rlabel polysilicon 14 5 14 5 3 A
rlabel ntransistor 14 7 14 7 3 A
rlabel polysilicon 14 17 14 17 3 A
rlabel ptransistor 14 24 14 24 3 A
rlabel polysilicon 14 54 14 54 3 A
rlabel ndiffusion 9 7 9 7 3 GND
rlabel pdiffusion 9 24 9 24 3 Vdd
rlabel m1 24 13 24 13 3 GND
rlabel m1 27 27 27 27 3 Y
port 1 e
rlabel m1 28 59 28 59 3 B
port 2 e
rlabel pdc 24 27 24 27 3 Y
port 1 e
rlabel pc 25 59 25 59 3 B
port 2 e
rlabel m1 25 63 25 63 3 B
port 2 e
rlabel m1 27 9 27 9 3 GND
rlabel m1 23 23 23 23 3 Y
port 1 e
rlabel m1 23 27 23 27 3 Y
port 1 e
rlabel m1 23 33 23 33 3 Y
port 1 e
rlabel m1 24 58 24 58 3 B
port 2 e
rlabel m1 24 59 24 59 3 B
port 2 e
rlabel m1 24 62 24 62 3 B
port 2 e
rlabel ndc 24 9 24 9 3 GND
rlabel m1 20 13 20 13 3 Y
port 1 e
rlabel m1 33 22 33 22 3 Y
port 1 e
rlabel ndc 17 13 17 13 3 Y
port 1 e
rlabel m1 17 47 17 47 3 Vdd
rlabel m1 16 12 16 12 3 Y
port 1 e
rlabel m1 16 13 16 13 3 Y
port 1 e
rlabel m1 16 16 16 16 3 Y
port 1 e
rlabel m1 16 18 16 18 3 Y
port 1 e
rlabel m1 16 22 16 22 3 Y
port 1 e
rlabel m1 13 44 13 44 3 Vdd
rlabel m1 13 47 13 47 3 Vdd
rlabel m1 13 59 13 59 3 A
port 3 e
rlabel ndc 10 9 10 9 3 GND
rlabel pdc 10 44 10 44 3 Vdd
rlabel pc 10 59 10 59 3 A
port 3 e
rlabel m1 9 5 9 5 3 GND
rlabel m1 9 9 9 9 3 GND
rlabel m1 9 13 9 13 3 GND
rlabel m1 9 43 9 43 3 Vdd
rlabel m1 9 44 9 44 3 Vdd
rlabel m1 9 49 9 49 3 Vdd
rlabel m1 9 58 9 58 3 A
port 3 e
rlabel m1 9 59 9 59 3 A
port 3 e
rlabel m1 9 62 9 62 3 A
port 3 e
rlabel m1 9 63 9 63 3 A
port 3 e
<< end >>
