VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005000 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 0.540000 BY 0.900000 ;
END CoreSite

LAYER m1
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.270000 ;
   WIDTH 0.270000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.270000 ;
   PITCH 0.540000 0.540000 ;
END m1

LAYER v1
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v1

LAYER m2
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m2

LAYER v2
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v2

LAYER m3
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m3

LAYER v3
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v3

LAYER m4
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m4

LAYER v4
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v4

LAYER m5
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m5

LAYER v5
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v5

LAYER m6
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m6

LAYER OVERLAP
   TYPE OVERLAP ;
END OVERLAP

VIA v1_C DEFAULT
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_C

VIA v1_Ch
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_Ch

VIA v1_Cv
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_Cv

VIA v2_C DEFAULT
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_C

VIA v2_Ch
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Ch

VIA v2_Cv
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Cv

VIA v3_C DEFAULT
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_C

VIA v3_Ch
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_Ch

VIA v3_Cv
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_Cv

VIA v4_C DEFAULT
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_C

VIA v4_Ch
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_Ch

VIA v4_Cv
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_Cv

VIA v5_C DEFAULT
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_C

VIA v5_Ch
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_Ch

VIA v5_Cv
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_Cv

MACRO _0_0cell_0_0g0n1n2naa_012aax0
    CLASS CORE ;
    FOREIGN _0_0cell_0_0g0n1n2naa_012aax0 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 7.020000 BY 8.100000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN in_50_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 6.570000 0.810000 7.740000 ;
        RECT 0.540000 6.480000 0.900000 6.570000 ;
        RECT 0.540000 6.300000 0.630000 6.480000 ;
        RECT 0.540000 6.210000 0.900000 6.300000 ;
        RECT 0.630000 6.300000 0.810000 6.480000 ;
        RECT 0.810000 6.300000 0.900000 6.480000 ;
        END
        ANTENNAGATEAREA 0.534600 ;
    END in_50_6
    PIN in_51_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 1.620000 7.020000 1.890000 7.740000 ;
        RECT 1.620000 6.930000 1.980000 7.020000 ;
        RECT 1.620000 6.750000 1.710000 6.930000 ;
        RECT 1.620000 6.660000 1.980000 6.750000 ;
        RECT 1.710000 6.750000 1.890000 6.930000 ;
        RECT 1.890000 6.750000 1.980000 6.930000 ;
        END
        ANTENNAGATEAREA 0.534600 ;
    END in_51_6
    PIN in_52_6
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 3.240000 6.660000 3.510000 7.740000 ;
        RECT 3.240000 6.570000 4.950000 6.660000 ;
        RECT 3.240000 6.390000 4.680000 6.570000 ;
        RECT 4.680000 6.390000 4.860000 6.570000 ;
        RECT 4.860000 6.390000 4.950000 6.570000 ;
        RECT 4.590000 6.300000 4.950000 6.390000 ;
        END
        ANTENNAGATEAREA 0.534600 ;
    END in_52_6
    PIN out
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.270000 1.890000 3.240000 2.070000 ;
        RECT 0.270000 1.800000 3.510000 1.890000 ;
        RECT 0.270000 1.530000 0.810000 1.800000 ;
        RECT 3.240000 1.890000 3.420000 2.070000 ;
        RECT 0.450000 0.810000 0.900000 1.170000 ;
        RECT 3.420000 1.890000 5.400000 2.070000 ;
        RECT 5.310000 1.800000 5.400000 1.890000 ;
        RECT 0.540000 1.170000 0.810000 1.530000 ;
        RECT 5.400000 1.800000 5.670000 2.070000 ;
        RECT 3.150000 2.070000 5.760000 2.160000 ;
        RECT 5.670000 1.800000 5.760000 2.070000 ;
        RECT 3.240000 2.160000 3.510000 4.320000 ;
        RECT 5.310000 1.710000 5.760000 1.800000 ;
        RECT 3.150000 4.590000 3.510000 4.680000 ;
        RECT 3.150000 4.410000 3.240000 4.590000 ;
        RECT 3.150000 4.320000 3.510000 4.410000 ;
        RECT 3.240000 4.410000 3.420000 4.590000 ;
        RECT 3.420000 4.410000 3.510000 4.590000 ;
        END
        ANTENNAGATEAREA 0.388800 ;
        ANTENNADIFFAREA 1.263600 ;
    END out
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.540000 4.590000 0.900000 4.680000 ;
        RECT 0.540000 4.410000 0.630000 4.590000 ;
        RECT 0.540000 4.320000 0.900000 4.410000 ;
        RECT 0.630000 5.580000 4.860000 5.760000 ;
        RECT 0.630000 5.490000 5.670000 5.580000 ;
        RECT 0.630000 4.680000 0.900000 5.490000 ;
        RECT 0.630000 4.410000 0.810000 4.590000 ;
        RECT 0.630000 3.510000 0.900000 4.320000 ;
        RECT 0.630000 3.420000 1.620000 3.510000 ;
        RECT 0.630000 3.240000 1.260000 3.420000 ;
        RECT 4.860000 5.580000 5.040000 5.760000 ;
        RECT 0.810000 4.410000 0.900000 4.590000 ;
        RECT 1.170000 3.150000 1.260000 3.240000 ;
        RECT 1.170000 3.060000 1.620000 3.150000 ;
        RECT 5.040000 5.580000 5.670000 5.760000 ;
        RECT 1.260000 3.150000 1.530000 3.420000 ;
        RECT 1.530000 3.150000 1.620000 3.420000 ;
        RECT 4.680000 5.850000 5.130000 5.940000 ;
        RECT 4.680000 5.760000 5.670000 5.850000 ;
        RECT 5.400000 5.850000 5.670000 7.740000 ;
        END
        ANTENNAGATEAREA 0.315900 ;
        ANTENNADIFFAREA 0.858600 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.540000 2.790000 0.900000 2.880000 ;
        RECT 0.540000 2.610000 0.630000 2.790000 ;
        RECT 0.540000 2.520000 2.610000 2.610000 ;
        RECT 0.630000 2.610000 0.810000 2.790000 ;
        RECT 2.610000 2.520000 2.880000 2.790000 ;
        RECT 0.810000 2.610000 2.610000 2.790000 ;
        RECT 2.880000 2.520000 2.970000 2.790000 ;
        RECT 2.520000 2.430000 2.970000 2.520000 ;
        RECT 1.170000 5.130000 1.620000 5.220000 ;
        RECT 1.170000 4.860000 1.260000 5.130000 ;
        RECT 1.170000 4.770000 2.160000 4.860000 ;
        RECT 1.260000 4.860000 1.530000 5.130000 ;
        RECT 1.530000 5.040000 1.620000 5.130000 ;
        RECT 1.530000 4.860000 2.160000 5.040000 ;
        RECT 1.890000 2.790000 2.160000 4.770000 ;
        RECT 6.300000 2.430000 6.750000 2.520000 ;
        RECT 4.680000 2.790000 5.130000 2.880000 ;
        RECT 4.680000 2.520000 4.770000 2.790000 ;
        RECT 4.680000 2.430000 5.130000 2.520000 ;
        RECT 2.520000 2.790000 2.970000 2.880000 ;
        RECT 4.770000 2.610000 4.860000 2.790000 ;
        RECT 4.770000 2.520000 5.040000 2.610000 ;
        RECT 4.860000 2.610000 5.040000 2.790000 ;
        RECT 5.040000 2.520000 5.130000 2.790000 ;
        RECT 6.300000 2.790000 6.750000 2.880000 ;
        RECT 6.300000 2.520000 6.390000 2.790000 ;
        RECT 6.480000 2.880000 6.750000 3.420000 ;
        RECT 6.390000 2.520000 6.660000 2.790000 ;
        RECT 6.660000 2.520000 6.750000 2.790000 ;
        LAYER v1 ;
        RECT 2.610000 2.520000 2.880000 2.790000 ;
        RECT 4.770000 2.610000 4.860000 2.790000 ;
        RECT 4.770000 2.520000 5.040000 2.610000 ;
        RECT 4.860000 2.610000 5.040000 2.790000 ;
        RECT 6.390000 2.520000 6.660000 2.790000 ;
        LAYER m2 ;
        RECT 2.520000 2.790000 6.750000 2.880000 ;
        RECT 2.520000 2.520000 2.610000 2.790000 ;
        RECT 2.520000 2.430000 6.750000 2.520000 ;
        RECT 2.610000 2.520000 2.880000 2.790000 ;
        RECT 2.880000 2.520000 4.770000 2.790000 ;
        RECT 4.770000 2.610000 4.860000 2.790000 ;
        RECT 4.770000 2.520000 5.040000 2.610000 ;
        RECT 4.860000 2.610000 5.040000 2.790000 ;
        RECT 5.040000 2.520000 6.390000 2.790000 ;
        RECT 6.390000 2.520000 6.660000 2.790000 ;
        RECT 6.660000 2.520000 6.750000 2.790000 ;
        END
        ANTENNAGATEAREA 0.145800 ;
        ANTENNADIFFAREA 0.761400 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 2.520000 5.130000 6.030000 5.220000 ;
        RECT 2.520000 4.950000 2.610000 5.130000 ;
        RECT 2.520000 4.860000 2.880000 4.950000 ;
        RECT 2.610000 4.950000 2.790000 5.130000 ;
        RECT 5.670000 4.590000 6.030000 4.680000 ;
        RECT 5.670000 4.410000 5.760000 4.590000 ;
        RECT 5.670000 4.320000 6.030000 4.410000 ;
        RECT 5.670000 2.880000 5.940000 4.320000 ;
        RECT 5.670000 2.790000 6.030000 2.880000 ;
        RECT 5.670000 2.520000 6.030000 2.610000 ;
        RECT 2.790000 4.950000 6.030000 5.130000 ;
        RECT 5.760000 4.680000 6.030000 4.950000 ;
        RECT 5.760000 4.410000 5.940000 4.590000 ;
        RECT 5.940000 4.410000 6.030000 4.590000 ;
        RECT 5.670000 2.610000 5.760000 2.790000 ;
        RECT 5.760000 2.610000 5.940000 2.790000 ;
        RECT 5.940000 2.610000 6.030000 2.790000 ;
    END
END _0_0cell_0_0g0n1n2naa_012aax0

MACRO welltap_svt
    CLASS CORE WELLTAP ;
    FOREIGN welltap_svt 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.620000 BY 2.700000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.540000 1.530000 0.810000 1.710000 ;
        RECT 0.540000 1.350000 0.990000 1.530000 ;
        RECT 0.540000 1.170000 0.630000 1.350000 ;
        RECT 0.540000 1.080000 0.990000 1.170000 ;
        RECT 0.810000 1.170000 0.990000 1.350000 ;
        END
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.540000 0.990000 0.630000 ;
        RECT 0.540000 0.270000 0.630000 0.540000 ;
        RECT 0.540000 0.180000 0.990000 0.270000 ;
        RECT 0.900000 0.270000 0.990000 0.540000 ;
        END
    END GND
END welltap_svt

MACRO circuitppnp
   CLASS CORE ;
   FOREIGN circuitppnp 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 244.620000 BY 259.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitppnp

MACRO circuitwell
   CLASS CORE ;
   FOREIGN circuitwell 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 244.620000 BY 259.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitwell

