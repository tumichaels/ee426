magic
tech TSMC180
timestamp 1734123549
<< ppdiff >>
rect 6 7 11 8
rect 6 4 7 7
rect 10 4 11 7
rect 6 3 11 4
<< nndiff >>
rect 6 16 11 18
rect 6 14 7 16
rect 9 14 11 16
rect 6 13 11 14
<< psubstratepcontact >>
rect 7 4 10 7
<< nsubstratencontact >>
rect 7 14 9 16
<< m1 >>
rect 6 18 9 20
rect 6 16 11 18
rect 6 14 7 16
rect 9 14 11 16
rect 6 13 11 14
rect 6 7 11 8
rect 6 4 7 7
rect 10 4 11 7
rect 6 3 11 4
<< labels >>
rlabel m1 7 18 7 18 3 Vdd
port 2 e
rlabel nndiff 7 14 7 14 3 Vdd
rlabel m1 6 3 7 8 2 GND
<< end >>
