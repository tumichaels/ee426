magic
tech sky130l
timestamp 1726537171
<< ndiffusion >>
rect 66 77 78 80
rect 66 71 69 77
rect 75 71 78 77
rect 66 68 78 71
rect 66 60 78 63
rect 66 54 69 60
rect 75 54 78 60
rect 66 51 78 54
<< ndc >>
rect 69 71 75 77
rect 69 54 75 60
<< ntransistor >>
rect 66 63 78 68
<< pdiffusion >>
rect 42 77 54 80
rect 42 71 45 77
rect 51 71 54 77
rect 42 68 54 71
rect 42 60 54 63
rect 42 54 45 60
rect 51 54 54 60
rect 42 51 54 54
<< pdc >>
rect 45 71 51 77
rect 45 54 51 60
<< ptransistor >>
rect 42 63 54 68
<< polysilicon >>
rect 40 63 42 68
rect 54 63 66 68
rect 78 63 86 68
<< m1 >>
rect 28 77 52 78
rect 28 71 45 77
rect 51 71 52 77
rect 28 70 52 71
rect 68 77 92 78
rect 68 71 69 77
rect 75 71 92 77
rect 68 70 92 71
rect 44 60 76 61
rect 44 54 45 60
rect 51 54 69 60
rect 75 54 76 60
rect 44 53 76 54
<< labels >>
rlabel m1 51 53 69 61 0 out
rlabel m1 28 70 45 78 1 Vdd!
rlabel m1 75 70 92 78 1 GND!
rlabel polysilicon 54 63 66 68 1 in
<< end >>
