magic
tech sky130l
timestamp 1731040975
<< ndiffusion >>
rect 8 14 13 16
rect 8 11 9 14
rect 12 11 13 14
rect 8 6 13 11
rect 15 6 20 16
rect 22 10 27 16
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 33 15 38 16
rect 33 12 34 15
rect 37 12 38 15
rect 33 6 38 12
rect 40 10 45 16
rect 40 7 41 10
rect 44 7 45 10
rect 40 6 45 7
rect 47 10 52 16
rect 47 7 48 10
rect 51 7 52 10
rect 47 6 52 7
rect 58 10 63 16
rect 58 7 59 10
rect 62 7 63 10
rect 58 6 63 7
rect 65 15 70 16
rect 65 12 66 15
rect 69 12 70 15
rect 65 6 70 12
<< ndc >>
rect 9 11 12 14
rect 23 7 26 10
rect 34 12 37 15
rect 41 7 44 10
rect 48 7 51 10
rect 59 7 62 10
rect 66 12 69 15
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 38 6 40 16
rect 45 6 47 16
rect 63 6 65 16
<< pdiffusion >>
rect 8 37 13 43
rect 8 34 9 37
rect 12 34 13 37
rect 8 23 13 34
rect 15 38 19 43
rect 15 37 20 38
rect 15 34 16 37
rect 19 34 20 37
rect 15 23 20 34
rect 22 27 27 38
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 33 27 38 33
rect 33 24 34 27
rect 37 24 38 27
rect 33 23 38 24
rect 40 23 45 33
rect 47 32 52 33
rect 47 29 48 32
rect 51 29 52 32
rect 47 23 52 29
rect 58 31 63 43
rect 58 28 59 31
rect 62 28 63 31
rect 58 23 63 28
rect 65 27 70 43
rect 65 24 66 27
rect 69 24 70 27
rect 65 23 70 24
<< pdc >>
rect 9 34 12 37
rect 16 34 19 37
rect 23 24 26 27
rect 34 24 37 27
rect 48 29 51 32
rect 59 28 62 31
rect 66 24 69 27
<< ptransistor >>
rect 13 23 15 43
rect 20 23 22 38
rect 38 23 40 33
rect 45 23 47 33
rect 63 23 65 43
<< polysilicon >>
rect 11 50 16 51
rect 11 47 12 50
rect 15 47 16 50
rect 11 46 16 47
rect 23 46 28 51
rect 65 50 70 51
rect 65 48 66 50
rect 63 47 66 48
rect 69 47 70 50
rect 13 43 15 46
rect 23 44 24 46
rect 20 43 24 44
rect 27 43 28 46
rect 20 42 28 43
rect 43 46 48 47
rect 43 43 44 46
rect 47 43 48 46
rect 63 46 70 47
rect 63 43 65 46
rect 43 42 48 43
rect 20 38 22 42
rect 38 33 40 35
rect 45 33 47 42
rect 13 16 15 23
rect 20 20 22 23
rect 38 20 40 23
rect 20 18 40 20
rect 20 16 22 18
rect 38 16 40 18
rect 45 16 47 23
rect 63 16 65 23
rect 13 4 15 6
rect 20 4 22 6
rect 38 4 40 6
rect 45 4 47 6
rect 63 4 65 6
<< pc >>
rect 12 47 15 50
rect 66 47 69 50
rect 24 43 27 46
rect 44 43 47 46
<< m1 >>
rect 11 50 16 51
rect 11 49 12 50
rect 8 47 12 49
rect 15 47 16 50
rect 8 46 16 47
rect 23 46 28 51
rect 8 44 12 46
rect 23 43 24 46
rect 27 43 28 46
rect 40 47 44 51
rect 66 50 69 51
rect 40 46 46 47
rect 40 44 44 46
rect 43 43 44 44
rect 47 43 48 46
rect 56 44 60 48
rect 66 46 69 47
rect 23 42 28 43
rect 9 37 12 38
rect 56 37 59 44
rect 15 34 16 37
rect 19 34 59 37
rect 9 33 12 34
rect 48 32 51 34
rect 48 28 51 29
rect 58 28 59 31
rect 62 28 63 31
rect 23 27 26 28
rect 66 27 69 28
rect 33 24 34 27
rect 37 24 38 27
rect 23 21 26 24
rect 23 18 37 21
rect 34 15 37 18
rect 66 15 69 24
rect 9 14 12 15
rect 33 12 34 15
rect 37 12 38 15
rect 66 11 69 12
rect 9 8 12 11
rect 8 4 12 8
rect 23 10 26 11
rect 41 10 44 11
rect 48 10 51 11
rect 26 7 41 9
rect 23 6 41 7
rect 44 6 45 9
rect 51 7 59 10
rect 62 7 63 10
rect 48 6 51 7
rect 40 5 45 6
rect 40 4 44 5
<< m2c >>
rect 66 47 69 50
rect 9 34 12 37
rect 59 28 62 31
rect 23 24 26 27
rect 34 24 37 27
rect 9 11 12 14
rect 66 12 69 15
rect 41 7 44 9
rect 41 6 44 7
<< m2 >>
rect 65 50 70 51
rect 65 47 66 50
rect 69 47 70 50
rect 65 46 70 47
rect 8 37 13 38
rect 8 34 9 37
rect 12 36 13 37
rect 12 34 60 36
rect 8 33 13 34
rect 58 32 60 34
rect 23 30 51 32
rect 23 28 25 30
rect 22 27 27 28
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 33 27 38 28
rect 33 24 34 27
rect 37 24 38 27
rect 33 23 38 24
rect 49 25 51 30
rect 58 31 63 32
rect 58 28 59 31
rect 62 28 63 31
rect 58 27 63 28
rect 66 25 68 46
rect 49 23 68 25
rect 35 15 37 23
rect 65 15 70 16
rect 8 14 66 15
rect 8 11 9 14
rect 12 13 66 14
rect 12 11 13 13
rect 65 12 66 13
rect 69 12 70 15
rect 65 11 70 12
rect 8 10 13 11
rect 40 9 45 10
rect 40 6 41 9
rect 44 6 45 9
rect 40 5 45 6
<< labels >>
rlabel space 0 0 80 56 6 prboundary
rlabel pdiffusion 70 25 70 25 3 _q
rlabel ndiffusion 66 7 66 7 3 _q
rlabel ndiffusion 59 8 59 8 3 #10
rlabel pdiffusion 66 24 66 24 3 _q
rlabel pdiffusion 66 25 66 25 3 _q
rlabel pdiffusion 66 28 66 28 3 _q
rlabel polysilicon 66 49 66 49 3 _clk
rlabel ntransistor 64 7 64 7 3 _clk
rlabel polysilicon 64 17 64 17 3 _clk
rlabel ptransistor 64 24 64 24 3 _clk
rlabel polysilicon 64 44 64 44 3 _clk
rlabel polysilicon 64 47 64 47 3 _clk
rlabel polysilicon 64 48 64 48 3 _clk
rlabel ndiffusion 59 7 59 7 3 #10
rlabel ndiffusion 59 11 59 11 3 #10
rlabel pdiffusion 59 24 59 24 3 #7
rlabel pdiffusion 52 30 52 30 3 Vdd
rlabel ndiffusion 48 7 48 7 3 #10
rlabel ndiffusion 48 8 48 8 3 #10
rlabel ndiffusion 48 11 48 11 3 #10
rlabel ndiffusion 45 8 45 8 3 GND
rlabel pdiffusion 48 24 48 24 3 Vdd
rlabel pdiffusion 48 30 48 30 3 Vdd
rlabel pdiffusion 48 33 48 33 3 Vdd
rlabel polysilicon 46 34 46 34 3 q
rlabel polysilicon 64 5 64 5 3 _clk
rlabel ntransistor 46 7 46 7 3 q
rlabel polysilicon 46 17 46 17 3 q
rlabel ptransistor 46 24 46 24 3 q
rlabel polysilicon 44 43 44 43 3 q
rlabel polysilicon 44 47 44 47 3 q
rlabel ndiffusion 41 8 41 8 3 GND
rlabel ndiffusion 41 11 41 11 3 GND
rlabel polysilicon 46 5 46 5 3 q
rlabel ntransistor 39 7 39 7 3 CLK
rlabel polysilicon 39 17 39 17 3 CLK
rlabel polysilicon 39 21 39 21 3 CLK
rlabel ptransistor 39 24 39 24 3 CLK
rlabel polysilicon 39 34 39 34 3 CLK
rlabel ndiffusion 34 7 34 7 3 _clk
rlabel ndiffusion 34 16 34 16 3 _clk
rlabel polysilicon 24 45 24 45 3 CLK
rlabel polysilicon 39 5 39 5 3 CLK
rlabel ndiffusion 23 7 23 7 3 GND
rlabel ndiffusion 23 8 23 8 3 GND
rlabel ndiffusion 23 11 23 11 3 GND
rlabel polysilicon 21 39 21 39 3 CLK
rlabel polysilicon 21 43 21 43 3 CLK
rlabel polysilicon 21 44 21 44 3 CLK
rlabel polysilicon 21 5 21 5 3 CLK
rlabel ntransistor 21 7 21 7 3 CLK
rlabel polysilicon 21 17 21 17 3 CLK
rlabel polysilicon 21 19 21 19 3 CLK
rlabel polysilicon 21 21 21 21 3 CLK
rlabel ptransistor 21 24 21 24 3 CLK
rlabel pdiffusion 16 24 16 24 3 Vdd
rlabel pdiffusion 16 38 16 38 3 Vdd
rlabel pdiffusion 16 39 16 39 3 Vdd
rlabel polysilicon 14 44 14 44 3 D
rlabel polysilicon 14 5 14 5 3 D
rlabel ntransistor 14 7 14 7 3 D
rlabel polysilicon 14 17 14 17 3 D
rlabel ptransistor 14 24 14 24 3 D
rlabel polysilicon 12 47 12 47 3 D
rlabel polysilicon 12 48 12 48 3 D
rlabel ndiffusion 9 7 9 7 3 _q
rlabel pdiffusion 9 24 9 24 3 #7
rlabel m1 67 47 67 47 3 _clk
rlabel m1 67 51 67 51 3 _clk
rlabel m1 67 16 67 16 3 _q
port 1 e
rlabel pdc 67 25 67 25 3 _q
port 1 e
rlabel m1 67 28 67 28 3 _q
port 1 e
rlabel m1 57 38 57 38 3 Vdd
rlabel m1 57 45 57 45 3 Vdd
rlabel m1 49 29 49 29 3 Vdd
rlabel pdc 49 30 49 30 3 Vdd
rlabel m1 49 33 49 33 3 Vdd
rlabel m1 48 44 48 44 3 q
port 2 e
rlabel pc 45 44 45 44 3 q
port 2 e
rlabel m1 44 44 44 44 3 q
port 2 e
rlabel m1 41 45 41 45 3 q
port 2 e
rlabel m1 41 47 41 47 3 q
port 2 e
rlabel m1 41 48 41 48 3 q
port 2 e
rlabel m1 63 8 63 8 3 #10
rlabel ndc 60 8 60 8 3 #10
rlabel m1 67 12 67 12 3 _q
port 1 e
rlabel m1 38 13 38 13 3 _clk
rlabel m1 28 44 28 44 3 CLK
port 3 e
rlabel m1 52 8 52 8 3 #10
rlabel ndc 35 13 35 13 3 _clk
rlabel m1 35 16 35 16 3 _clk
rlabel pc 25 44 25 44 3 CLK
port 3 e
rlabel m1 49 7 49 7 3 #10
rlabel ndc 49 8 49 8 3 #10
rlabel m1 49 11 49 11 3 #10
rlabel m1 34 13 34 13 3 _clk
rlabel m1 24 43 24 43 3 CLK
port 3 e
rlabel m1 24 44 24 44 3 CLK
port 3 e
rlabel m1 24 47 24 47 3 CLK
port 3 e
rlabel m1 24 19 24 19 3 _clk
rlabel m1 24 22 24 22 3 _clk
rlabel m1 24 28 24 28 3 _clk
rlabel m1 20 35 20 35 3 Vdd
rlabel ndc 42 10 42 10 3 GND
rlabel m1 42 11 42 11 3 GND
rlabel pdc 17 35 17 35 3 Vdd
rlabel m1 41 5 41 5 3 GND
rlabel m1 27 8 27 8 3 GND
rlabel m1 24 11 24 11 3 GND
rlabel m1 16 35 16 35 3 Vdd
rlabel m1 24 7 24 7 3 GND
rlabel ndc 24 8 24 8 3 GND
rlabel m1 16 48 16 48 3 D
port 4 e
rlabel m1 12 50 12 50 3 D
port 4 e
rlabel m1 12 51 12 51 3 D
port 4 e
rlabel m1 10 9 10 9 3 _q
port 1 e
rlabel m1 10 15 10 15 3 _q
port 1 e
rlabel m1 10 34 10 34 3 #7
rlabel m1 10 38 10 38 3 #7
rlabel pc 13 48 13 48 3 D
port 4 e
rlabel m1 9 5 9 5 3 _q
port 1 e
rlabel m1 9 45 9 45 3 D
port 4 e
rlabel m1 9 47 9 47 3 D
port 4 e
rlabel m1 9 48 9 48 3 D
port 4 e
rlabel m2 67 26 67 26 3 _clk
rlabel m2 63 29 63 29 3 #7
rlabel m2c 60 29 60 29 3 #7
rlabel m2 59 28 59 28 3 #7
rlabel m2 59 29 59 29 3 #7
rlabel m2 66 16 66 16 3 _q
port 1 e
rlabel m2 50 26 50 26 3 _clk
rlabel m2 70 13 70 13 3 _q
port 1 e
rlabel m2 50 24 50 24 3 _clk
rlabel m2 38 25 38 25 3 _q
port 1 e
rlabel m2c 67 13 67 13 3 _q
port 1 e
rlabel m2c 35 25 35 25 3 _q
port 1 e
rlabel m2 66 12 66 12 3 _q
port 1 e
rlabel m2 66 13 66 13 3 _q
port 1 e
rlabel m2 34 25 34 25 3 _q
port 1 e
rlabel m2 45 7 45 7 3 GND
rlabel m2 59 32 59 32 3 #7
rlabel m2 59 33 59 33 3 #7
rlabel m2c 42 7 42 7 3 GND
rlabel m2c 42 8 42 8 3 GND
rlabel m2 36 16 36 16 3 _q
port 1 e
rlabel m2 34 24 34 24 3 _q
port 1 e
rlabel m2 27 25 27 25 3 _clk
rlabel m2 34 28 34 28 3 _q
port 1 e
rlabel m2 41 6 41 6 3 GND
rlabel m2 41 7 41 7 3 GND
rlabel m2 41 10 41 10 3 GND
rlabel m2c 24 25 24 25 3 _clk
rlabel m2 24 29 24 29 3 _clk
rlabel m2 24 31 24 31 3 _clk
rlabel m2 70 48 70 48 3 _clk
rlabel m2 23 24 23 24 3 _clk
rlabel m2 23 25 23 25 3 _clk
rlabel m2 23 28 23 28 3 _clk
rlabel m2c 67 48 67 48 3 _clk
rlabel m2 13 12 13 12 3 _q
port 1 e
rlabel m2 13 14 13 14 3 _q
port 1 e
rlabel m2 13 35 13 35 3 #7
rlabel m2 13 37 13 37 3 #7
rlabel m2 66 47 66 47 3 _clk
rlabel m2 66 48 66 48 3 _clk
rlabel m2 66 51 66 51 3 _clk
rlabel m2c 10 12 10 12 3 _q
port 1 e
rlabel m2c 10 35 10 35 3 #7
rlabel m2 9 11 9 11 3 _q
port 1 e
rlabel m2 9 12 9 12 3 _q
port 1 e
rlabel m2 9 15 9 15 3 _q
port 1 e
rlabel m2 9 34 9 34 3 #7
rlabel m2 9 35 9 35 3 #7
rlabel m2 9 38 9 38 3 #7
<< end >>
