VERSION 5.6 ;

BUSBITCHARS "[]" ;

DIVIDERCHAR "/" ;

UNITS
    DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005000 ; 

CLEARANCEMEASURE EUCLIDEAN ; 

USEMINSPACING OBS ON ; 

SITE CoreSite
    CLASS CORE ;
    SIZE 0.540000 BY 0.900000 ;
END CoreSite

LAYER m1
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.270000 ;
   WIDTH 0.270000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.270000 ;
   PITCH 0.540000 0.540000 ;
END m1

LAYER v1
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v1

LAYER m2
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m2

LAYER v2
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v2

LAYER m3
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m3

LAYER v3
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v3

LAYER m4
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m4

LAYER v4
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v4

LAYER m5
   TYPE ROUTING ;
   DIRECTION VERTICAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m5

LAYER v5
    TYPE CUT ;
    SPACING 0.270000 ;
    WIDTH 0.270000 ;
    ENCLOSURE ABOVE 0.090000 0.090000 ;
    ENCLOSURE BELOW 0.090000 0.090000 ;
END v5

LAYER m6
   TYPE ROUTING ;
   DIRECTION HORIZONTAL ;
   MINWIDTH 0.450000 ;
   WIDTH 0.450000 ;
   SPACINGTABLE
      PARALLELRUNLENGTH 0.0
      WIDTH 0.0 0.450000 ;
   PITCH 0.900000 0.900000 ;
END m6

LAYER OVERLAP
   TYPE OVERLAP ;
END OVERLAP

VIA v1_C DEFAULT
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_C

VIA v1_Ch
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_Ch

VIA v1_Cv
   LAYER m1 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v1 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v1_Cv

VIA v2_C DEFAULT
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_C

VIA v2_Ch
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Ch

VIA v2_Cv
   LAYER m2 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v2 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v2_Cv

VIA v3_C DEFAULT
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_C

VIA v3_Ch
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_Ch

VIA v3_Cv
   LAYER m3 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v3 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v3_Cv

VIA v4_C DEFAULT
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_C

VIA v4_Ch
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_Ch

VIA v4_Cv
   LAYER m4 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v4 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v4_Cv

VIA v5_C DEFAULT
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_C

VIA v5_Ch
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_Ch

VIA v5_Cv
   LAYER m5 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
   LAYER v5 ;
     RECT -0.135000 -0.135000 0.135000 0.135000 ;
   LAYER m6 ;
     RECT -0.225000 -0.225000 0.225000 0.225000 ;
END v5_Cv

MACRO _0_0std_0_0cells_0_0AND2X1
    CLASS CORE ;
    FOREIGN _0_0std_0_0cells_0_0AND2X1 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 4.320000 BY 7.200000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN A
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 0.540000 6.030000 0.810000 6.300000 ;
        RECT 0.540000 5.940000 0.900000 6.030000 ;
        RECT 0.540000 5.760000 0.630000 5.940000 ;
        RECT 0.540000 5.670000 0.900000 5.760000 ;
        RECT 0.630000 5.760000 0.810000 5.940000 ;
        RECT 0.810000 5.760000 0.900000 5.940000 ;
        END
        ANTENNAGATEAREA 0.291600 ;
    END A
    PIN B
        DIRECTION INPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.610000 6.030000 2.970000 6.120000 ;
        RECT 2.610000 5.850000 2.700000 6.030000 ;
        RECT 2.610000 5.760000 2.970000 5.850000 ;
        RECT 2.700000 6.120000 2.970000 6.300000 ;
        RECT 2.700000 5.850000 2.880000 6.030000 ;
        RECT 2.880000 5.850000 2.970000 6.030000 ;
        END
        ANTENNAGATEAREA 0.291600 ;
    END B
    PIN Y
        DIRECTION OUTPUT ;
        USE SIGNAL ;
        PORT
        LAYER m1 ;
        RECT 2.700000 0.990000 2.970000 1.980000 ;
        RECT 2.700000 1.980000 3.060000 2.520000 ;
        RECT 2.700000 2.520000 2.790000 2.700000 ;
        RECT 2.790000 2.520000 2.970000 2.700000 ;
        RECT 2.970000 2.520000 3.060000 2.700000 ;
        RECT 2.700000 4.590000 3.060000 4.680000 ;
        RECT 2.700000 4.410000 2.790000 4.590000 ;
        RECT 2.700000 4.320000 3.060000 4.410000 ;
        RECT 2.700000 2.790000 2.970000 4.320000 ;
        RECT 2.700000 2.700000 3.060000 2.790000 ;
        RECT 2.790000 4.410000 2.970000 4.590000 ;
        RECT 2.970000 4.410000 3.060000 4.590000 ;
        END
        ANTENNADIFFAREA 0.631800 ;
    END Y
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.720000 4.950000 1.080000 5.040000 ;
        RECT 0.720000 4.770000 0.810000 4.950000 ;
        RECT 0.720000 4.680000 1.080000 4.770000 ;
        RECT 0.810000 5.130000 2.250000 5.400000 ;
        RECT 0.810000 5.040000 1.080000 5.130000 ;
        RECT 0.810000 4.770000 0.990000 4.950000 ;
        RECT 0.990000 4.770000 1.080000 4.950000 ;
        RECT 1.350000 5.760000 1.890000 6.030000 ;
        RECT 1.350000 5.400000 1.620000 5.760000 ;
        RECT 1.620000 6.030000 1.890000 6.300000 ;
        RECT 1.980000 5.040000 2.250000 5.130000 ;
        RECT 1.980000 4.950000 2.340000 5.040000 ;
        RECT 1.980000 4.770000 2.070000 4.950000 ;
        RECT 1.980000 4.680000 2.340000 4.770000 ;
        RECT 2.070000 4.770000 2.250000 4.950000 ;
        RECT 2.250000 4.770000 2.340000 4.950000 ;
        END
        ANTENNADIFFAREA 0.777600 ;
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 1.980000 2.520000 2.430000 2.610000 ;
        RECT 1.980000 2.880000 2.430000 2.970000 ;
        RECT 1.980000 2.610000 2.070000 2.880000 ;
        RECT 2.070000 2.790000 2.340000 2.880000 ;
        RECT 2.070000 2.610000 2.160000 2.790000 ;
        RECT 2.160000 2.610000 2.340000 2.790000 ;
        RECT 3.330000 2.610000 3.420000 2.880000 ;
        RECT 3.330000 2.520000 3.780000 2.610000 ;
        RECT 2.340000 2.610000 2.430000 2.880000 ;
        RECT 3.420000 2.610000 3.690000 2.880000 ;
        RECT 3.690000 2.610000 3.780000 2.880000 ;
        RECT 3.510000 6.030000 4.050000 6.300000 ;
        RECT 3.330000 2.880000 3.780000 2.970000 ;
        RECT 3.510000 2.970000 3.780000 6.030000 ;
        LAYER v1 ;
        RECT 2.070000 2.790000 2.340000 2.880000 ;
        RECT 2.070000 2.610000 2.160000 2.790000 ;
        RECT 2.160000 2.610000 2.340000 2.790000 ;
        RECT 3.420000 2.610000 3.690000 2.880000 ;
        LAYER m2 ;
        RECT 1.980000 2.880000 3.780000 2.970000 ;
        RECT 1.980000 2.610000 2.070000 2.880000 ;
        RECT 1.980000 2.520000 3.780000 2.610000 ;
        RECT 2.070000 2.790000 2.340000 2.880000 ;
        RECT 2.070000 2.610000 2.160000 2.790000 ;
        RECT 2.160000 2.610000 2.340000 2.790000 ;
        RECT 2.340000 2.610000 3.420000 2.880000 ;
        RECT 3.420000 2.610000 3.690000 2.880000 ;
        RECT 3.690000 2.610000 3.780000 2.880000 ;
        END
        ANTENNADIFFAREA 0.405000 ;
    END GND
    OBS
        LAYER m1 ;
        RECT 0.360000 1.350000 0.720000 1.440000 ;
        RECT 0.360000 1.170000 0.450000 1.350000 ;
        RECT 0.360000 1.080000 0.720000 1.170000 ;
        RECT 0.450000 1.440000 0.990000 1.710000 ;
        RECT 0.450000 1.170000 0.630000 1.350000 ;
        RECT 0.630000 1.170000 0.720000 1.350000 ;
        RECT 0.630000 1.710000 0.990000 1.800000 ;
        RECT 0.720000 2.790000 1.080000 2.880000 ;
        RECT 0.720000 2.610000 0.810000 2.790000 ;
        RECT 0.720000 2.520000 1.080000 2.610000 ;
        RECT 0.720000 1.800000 0.990000 2.520000 ;
        RECT 0.810000 4.140000 1.710000 4.410000 ;
        RECT 0.810000 2.880000 1.080000 4.140000 ;
        RECT 0.810000 2.610000 0.990000 2.790000 ;
        RECT 0.990000 2.610000 1.080000 2.790000 ;
        RECT 1.350000 4.590000 1.710000 4.680000 ;
        RECT 1.350000 4.410000 1.440000 4.590000 ;
        RECT 1.440000 4.410000 1.620000 4.590000 ;
        RECT 1.620000 4.410000 1.710000 4.590000 ;
    END
END _0_0std_0_0cells_0_0AND2X1

MACRO welltap_svt
    CLASS CORE WELLTAP ;
    FOREIGN welltap_svt 0.000000 0.000000 ;
    ORIGIN 0.000000 0.000000 ;
    SIZE 1.620000 BY 2.700000 ;
    SYMMETRY X Y ;
    SITE CoreSite ;
    PIN Vdd
        DIRECTION INPUT ;
        USE POWER ;
        PORT
        LAYER m1 ;
        RECT 0.540000 1.530000 0.810000 1.710000 ;
        RECT 0.540000 1.350000 0.990000 1.530000 ;
        RECT 0.540000 1.170000 0.630000 1.350000 ;
        RECT 0.540000 1.080000 0.990000 1.170000 ;
        RECT 0.810000 1.170000 0.990000 1.350000 ;
        END
    END Vdd
    PIN GND
        DIRECTION INPUT ;
        USE GROUND ;
        PORT
        LAYER m1 ;
        RECT 0.540000 0.540000 0.990000 0.630000 ;
        RECT 0.540000 0.270000 0.630000 0.540000 ;
        RECT 0.540000 0.180000 0.990000 0.270000 ;
        RECT 0.900000 0.270000 0.990000 0.540000 ;
        END
    END GND
END welltap_svt

MACRO circuitppnp
   CLASS CORE ;
   FOREIGN circuitppnp 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 255.960000 BY 259.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitppnp

MACRO circuitwell
   CLASS CORE ;
   FOREIGN circuitwell 0.000000 0.000000 ;
   ORIGIN 0.000000 0.000000 ; 
   SIZE 255.960000 BY 259.200000 ; 
   SYMMETRY X Y ;
   SITE CoreSite ;
END circuitwell

