magic
tech sky130l
timestamp 1731009265
<< ndiffusion >>
rect 8 10 13 16
rect 8 7 9 10
rect 12 7 13 10
rect 8 6 13 7
rect 15 6 20 16
rect 22 10 27 16
rect 22 7 23 10
rect 26 7 27 10
rect 22 6 27 7
rect 33 15 38 16
rect 33 12 34 15
rect 37 12 38 15
rect 33 6 38 12
rect 40 10 45 16
rect 40 7 41 10
rect 44 7 45 10
rect 40 6 45 7
rect 47 10 52 16
rect 47 7 48 10
rect 51 7 52 10
rect 47 6 52 7
rect 58 10 63 16
rect 58 7 59 10
rect 62 7 63 10
rect 58 6 63 7
rect 65 15 70 16
rect 65 12 66 15
rect 69 12 70 15
rect 65 6 70 12
<< ndc >>
rect 9 7 12 10
rect 23 7 26 10
rect 34 12 37 15
rect 41 7 44 10
rect 48 7 51 10
rect 59 7 62 10
rect 66 12 69 15
<< ntransistor >>
rect 13 6 15 16
rect 20 6 22 16
rect 38 6 40 16
rect 45 6 47 16
rect 63 6 65 16
<< pdiffusion >>
rect 8 28 13 43
rect 8 25 9 28
rect 12 25 13 28
rect 8 23 13 25
rect 15 38 19 43
rect 15 27 20 38
rect 15 24 16 27
rect 19 24 20 27
rect 15 23 20 24
rect 22 27 27 38
rect 22 24 23 27
rect 26 24 27 27
rect 22 23 27 24
rect 33 27 38 33
rect 33 24 34 27
rect 37 24 38 27
rect 33 23 38 24
rect 40 23 45 33
rect 47 32 52 33
rect 47 29 48 32
rect 51 29 52 32
rect 47 23 52 29
rect 58 27 63 43
rect 58 24 59 27
rect 62 24 63 27
rect 58 23 63 24
rect 65 40 70 43
rect 65 37 66 40
rect 69 37 70 40
rect 65 23 70 37
<< pdc >>
rect 9 25 12 28
rect 16 24 19 27
rect 23 24 26 27
rect 34 24 37 27
rect 48 29 51 32
rect 59 24 62 27
rect 66 37 69 40
<< ptransistor >>
rect 13 23 15 43
rect 20 23 22 38
rect 38 23 40 33
rect 45 23 47 33
rect 63 23 65 43
<< polysilicon >>
rect 24 47 29 48
rect 24 46 25 47
rect 13 44 25 46
rect 28 44 29 47
rect 13 43 15 44
rect 24 43 29 44
rect 40 47 45 48
rect 40 44 41 47
rect 44 44 45 47
rect 40 43 45 44
rect 48 47 53 48
rect 48 44 49 47
rect 52 45 53 47
rect 52 44 56 45
rect 48 43 56 44
rect 63 43 65 45
rect 32 40 37 41
rect 20 38 22 40
rect 32 37 33 40
rect 36 38 37 40
rect 36 37 40 38
rect 32 36 40 37
rect 38 33 40 36
rect 43 37 45 43
rect 43 35 47 37
rect 45 33 47 35
rect 13 16 15 23
rect 20 21 22 23
rect 38 21 40 23
rect 20 19 40 21
rect 20 16 22 19
rect 38 16 40 19
rect 45 16 47 23
rect 54 21 56 43
rect 63 21 65 23
rect 54 19 65 21
rect 63 16 65 19
rect 13 4 15 6
rect 20 4 22 6
rect 38 4 40 6
rect 45 4 47 6
rect 63 4 65 6
<< pc >>
rect 25 44 28 47
rect 41 44 44 47
rect 49 44 52 47
rect 33 37 36 40
<< m1 >>
rect 8 47 12 48
rect 8 44 9 47
rect 24 47 28 48
rect 40 47 44 48
rect 24 44 25 47
rect 28 44 29 47
rect 40 44 41 47
rect 41 43 44 44
rect 49 47 52 48
rect 56 47 60 48
rect 56 44 57 47
rect 72 44 76 48
rect 49 43 52 44
rect 33 40 36 41
rect 66 40 69 41
rect 33 36 36 37
rect 49 37 66 40
rect 49 32 52 37
rect 9 28 12 29
rect 9 21 12 25
rect 16 27 19 28
rect 16 23 19 24
rect 23 27 26 32
rect 47 29 48 32
rect 51 29 52 32
rect 23 16 26 24
rect 34 27 37 28
rect 34 23 37 24
rect 59 27 62 28
rect 59 23 62 24
rect 23 15 38 16
rect 23 13 34 15
rect 33 12 34 13
rect 37 12 38 15
rect 66 15 69 37
rect 66 11 69 12
rect 9 10 12 11
rect 41 10 44 11
rect 48 10 51 11
rect 59 10 62 11
rect 8 7 9 8
rect 8 4 12 7
rect 22 7 23 10
rect 26 9 28 10
rect 26 7 41 9
rect 44 7 45 10
rect 22 6 45 7
rect 51 7 59 10
rect 62 7 63 10
rect 48 6 51 7
rect 59 6 62 7
<< m2c >>
rect 9 44 12 47
rect 49 44 52 47
rect 57 44 60 47
rect 72 41 75 44
rect 33 37 36 40
rect 23 32 26 35
rect 16 24 19 27
rect 9 18 12 21
rect 34 24 37 27
rect 59 24 62 27
rect 41 7 44 10
<< m2 >>
rect 8 47 13 48
rect 48 47 53 48
rect 8 44 9 47
rect 12 45 34 47
rect 48 45 49 47
rect 12 44 13 45
rect 8 43 13 44
rect 32 41 34 45
rect 39 44 49 45
rect 52 44 53 47
rect 39 43 53 44
rect 56 47 61 48
rect 56 44 57 47
rect 60 44 61 47
rect 56 43 61 44
rect 71 44 76 45
rect 32 40 37 41
rect 32 37 33 40
rect 36 37 37 40
rect 32 36 37 37
rect 22 35 27 36
rect 22 32 23 35
rect 26 34 27 35
rect 39 34 41 43
rect 56 41 58 43
rect 26 32 41 34
rect 43 39 58 41
rect 71 41 72 44
rect 75 41 76 44
rect 71 40 76 41
rect 22 31 27 32
rect 43 30 45 39
rect 35 28 45 30
rect 15 27 38 28
rect 15 24 16 27
rect 19 26 34 27
rect 19 24 20 26
rect 15 23 20 24
rect 33 24 34 26
rect 37 24 38 27
rect 33 23 38 24
rect 58 27 63 28
rect 58 24 59 27
rect 62 24 63 27
rect 58 23 63 24
rect 8 21 13 22
rect 8 18 9 21
rect 12 20 13 21
rect 58 20 60 23
rect 12 18 60 20
rect 8 17 13 18
rect 40 10 45 11
rect 40 7 41 10
rect 44 8 45 10
rect 74 8 76 40
rect 44 7 76 8
rect 40 6 76 7
<< labels >>
rlabel space 0 0 80 52 6 prboundary
rlabel pdiffusion 70 38 70 38 3 _q
rlabel polysilicon 64 44 64 44 3 _clk
rlabel polysilicon 53 46 53 46 3 _clk
rlabel ndiffusion 70 13 70 13 3 _q
rlabel pdiffusion 66 24 66 24 3 _q
rlabel pdiffusion 66 38 66 38 3 _q
rlabel pdiffusion 66 41 66 41 3 _q
rlabel polysilicon 64 22 64 22 3 _clk
rlabel ptransistor 64 24 64 24 3 _clk
rlabel polysilicon 49 44 49 44 3 _clk
rlabel polysilicon 49 45 49 45 3 _clk
rlabel ndiffusion 66 7 66 7 3 _q
rlabel ndiffusion 66 13 66 13 3 _q
rlabel ndiffusion 66 16 66 16 3 _q
rlabel ndiffusion 59 8 59 8 3 #10
rlabel polysilicon 64 17 64 17 3 _clk
rlabel polysilicon 45 45 45 45 3 q
rlabel ntransistor 64 7 64 7 3 _clk
rlabel polysilicon 46 34 46 34 3 q
rlabel ndiffusion 59 7 59 7 3 #10
rlabel ndiffusion 59 11 59 11 3 #10
rlabel polysilicon 55 20 55 20 3 _clk
rlabel polysilicon 55 22 55 22 3 _clk
rlabel pdiffusion 48 24 48 24 3 _q
rlabel pdiffusion 48 33 48 33 3 _q
rlabel polysilicon 44 36 44 36 3 q
rlabel polysilicon 44 38 44 38 3 q
rlabel polysilicon 41 44 41 44 3 q
rlabel polysilicon 46 17 46 17 3 q
rlabel ptransistor 46 24 46 24 3 q
rlabel ndiffusion 48 7 48 7 3 #10
rlabel ndiffusion 48 8 48 8 3 #10
rlabel ndiffusion 48 11 48 11 3 #10
rlabel polysilicon 39 34 39 34 3 CLK
rlabel polysilicon 64 5 64 5 3 _clk
rlabel ntransistor 46 7 46 7 3 q
rlabel polysilicon 39 17 39 17 3 CLK
rlabel polysilicon 39 22 39 22 3 CLK
rlabel ptransistor 39 24 39 24 3 CLK
rlabel polysilicon 37 39 37 39 3 CLK
rlabel ndiffusion 34 16 34 16 3 _clk
rlabel pdiffusion 34 28 34 28 3 Vdd
rlabel polysilicon 46 5 46 5 3 q
rlabel ntransistor 39 7 39 7 3 CLK
rlabel ndiffusion 34 7 34 7 3 _clk
rlabel pdiffusion 27 25 27 25 3 _clk
rlabel polysilicon 25 44 25 44 3 D
rlabel polysilicon 25 47 25 47 3 D
rlabel polysilicon 39 5 39 5 3 CLK
rlabel ndiffusion 23 11 23 11 3 GND
rlabel pdiffusion 23 24 23 24 3 _clk
rlabel pdiffusion 23 25 23 25 3 _clk
rlabel pdiffusion 23 28 23 28 3 _clk
rlabel polysilicon 21 39 21 39 3 CLK
rlabel polysilicon 21 5 21 5 3 CLK
rlabel ntransistor 21 7 21 7 3 CLK
rlabel polysilicon 21 17 21 17 3 CLK
rlabel polysilicon 21 20 21 20 3 CLK
rlabel polysilicon 21 22 21 22 3 CLK
rlabel ptransistor 21 24 21 24 3 CLK
rlabel ndiffusion 13 8 13 8 3 _q
rlabel pdiffusion 16 39 16 39 3 Vdd
rlabel pdiffusion 13 26 13 26 3 #7
rlabel polysilicon 14 5 14 5 3 D
rlabel ntransistor 14 7 14 7 3 D
rlabel polysilicon 14 17 14 17 3 D
rlabel ptransistor 14 24 14 24 3 D
rlabel polysilicon 14 44 14 44 3 D
rlabel polysilicon 14 45 14 45 3 D
rlabel ndiffusion 9 7 9 7 3 _q
rlabel ndiffusion 9 11 9 11 3 _q
rlabel pdiffusion 9 24 9 24 3 #7
rlabel pdiffusion 9 26 9 26 3 #7
rlabel pdiffusion 9 29 9 29 3 #7
rlabel m1 73 45 73 45 3 GND
rlabel m1 67 41 67 41 3 _q
port 1 e
rlabel ndc 67 13 67 13 3 _q
port 1 e
rlabel m1 67 16 67 16 3 _q
port 1 e
rlabel pdc 67 38 67 38 3 _q
port 1 e
rlabel m1 60 24 60 24 3 #7
rlabel m1 60 28 60 28 3 #7
rlabel m1 52 30 52 30 3 _q
port 1 e
rlabel m1 50 33 50 33 3 _q
port 1 e
rlabel m1 50 38 50 38 3 _q
port 1 e
rlabel m1 50 44 50 44 3 _clk
rlabel m1 50 48 50 48 3 _clk
rlabel m1 67 12 67 12 3 _q
port 1 e
rlabel pdc 49 30 49 30 3 _q
port 1 e
rlabel m1 48 30 48 30 3 _q
port 1 e
rlabel m1 63 8 63 8 3 #10
rlabel m1 42 44 42 44 3 q
port 2 e
rlabel ndc 60 8 60 8 3 #10
rlabel m1 60 11 60 11 3 #10
rlabel m1 52 8 52 8 3 #10
rlabel ndc 49 8 49 8 3 #10
rlabel m1 49 11 49 11 3 #10
rlabel m1 42 11 42 11 3 GND
rlabel m1 38 13 38 13 3 _clk
rlabel ndc 35 13 35 13 3 _clk
rlabel m1 34 13 34 13 3 _clk
rlabel pc 42 45 42 45 3 q
port 2 e
rlabel m1 35 24 35 24 3 Vdd
rlabel m1 35 28 35 28 3 Vdd
rlabel m1 29 45 29 45 3 D
port 3 e
rlabel m1 41 45 41 45 3 q
port 2 e
rlabel m1 41 48 41 48 3 q
port 2 e
rlabel m1 34 37 34 37 3 CLK
port 4 e
rlabel m1 34 41 34 41 3 CLK
port 4 e
rlabel pc 26 45 26 45 3 D
port 3 e
rlabel m1 60 7 60 7 3 #10
rlabel m1 27 8 27 8 3 GND
rlabel m1 27 10 27 10 3 GND
rlabel m1 25 45 25 45 3 D
port 3 e
rlabel m1 25 48 25 48 3 D
port 3 e
rlabel ndc 24 8 24 8 3 GND
rlabel m1 24 14 24 14 3 _clk
rlabel m1 24 16 24 16 3 _clk
rlabel m1 24 17 24 17 3 _clk
rlabel pdc 24 25 24 25 3 _clk
rlabel m1 24 28 24 28 3 _clk
rlabel m1 49 7 49 7 3 #10
rlabel m1 23 8 23 8 3 GND
rlabel m1 17 24 17 24 3 Vdd
rlabel m1 17 28 17 28 3 Vdd
rlabel m1 23 7 23 7 3 GND
rlabel ndc 10 8 10 8 3 _q
port 1 e
rlabel m1 10 11 10 11 3 _q
port 1 e
rlabel m1 10 22 10 22 3 #7
rlabel pdc 10 26 10 26 3 #7
rlabel m1 10 29 10 29 3 #7
rlabel m1 9 5 9 5 3 _q
port 1 e
rlabel m1 9 8 9 8 3 _q
port 1 e
rlabel m2 76 42 76 42 3 GND
rlabel m2c 73 42 73 42 3 GND
rlabel m2 72 42 72 42 3 GND
rlabel m2 72 41 72 41 3 GND
rlabel m2 72 45 72 45 3 GND
rlabel m2 57 42 57 42 3 Vdd
rlabel m2 63 25 63 25 3 #7
rlabel m2 44 40 44 40 3 Vdd
rlabel m2 61 45 61 45 3 Vdd
rlabel m2c 60 25 60 25 3 #7
rlabel m2c 58 45 58 45 3 Vdd
rlabel m2 59 25 59 25 3 #7
rlabel m2 59 28 59 28 3 #7
rlabel m2 40 35 40 35 3 _clk
rlabel m2 57 45 57 45 3 Vdd
rlabel m2 75 9 75 9 3 GND
rlabel m2 44 31 44 31 3 Vdd
rlabel m2 59 21 59 21 3 #7
rlabel m2 59 24 59 24 3 #7
rlabel m2 57 44 57 44 3 Vdd
rlabel m2 53 45 53 45 3 _clk
rlabel m2c 50 45 50 45 3 _clk
rlabel m2 38 25 38 25 3 Vdd
rlabel m2 36 29 36 29 3 Vdd
rlabel m2 37 38 37 38 3 CLK
port 4 e
rlabel m2 40 44 40 44 3 _clk
rlabel m2 40 45 40 45 3 _clk
rlabel m2 45 8 45 8 3 GND
rlabel m2 45 9 45 9 3 GND
rlabel m2c 35 25 35 25 3 Vdd
rlabel m2c 34 38 34 38 3 CLK
port 4 e
rlabel m2c 42 8 42 8 3 GND
rlabel m2 34 24 34 24 3 Vdd
rlabel m2 34 25 34 25 3 Vdd
rlabel m2 27 33 27 33 3 _clk
rlabel m2 27 35 27 35 3 _clk
rlabel m2 33 37 33 37 3 CLK
port 4 e
rlabel m2 33 38 33 38 3 CLK
port 4 e
rlabel m2 33 41 33 41 3 CLK
port 4 e
rlabel m2 33 42 33 42 3 CLK
port 4 e
rlabel m2 41 7 41 7 3 GND
rlabel m2 41 8 41 8 3 GND
rlabel m2 41 11 41 11 3 GND
rlabel m2c 24 33 24 33 3 _clk
rlabel m2 23 32 23 32 3 _clk
rlabel m2 23 33 23 33 3 _clk
rlabel m2 23 36 23 36 3 _clk
rlabel m2 20 25 20 25 3 Vdd
rlabel m2 20 27 20 27 3 Vdd
rlabel m2 49 46 49 46 3 _clk
rlabel m2 57 48 57 48 3 Vdd
rlabel m2c 17 25 17 25 3 Vdd
rlabel m2 13 19 13 19 3 #7
rlabel m2 13 21 13 21 3 #7
rlabel m2 16 24 16 24 3 Vdd
rlabel m2 16 25 16 25 3 Vdd
rlabel m2 16 28 16 28 3 Vdd
rlabel m2 13 45 13 45 3 CLK
port 4 e
rlabel m2 13 46 13 46 3 CLK
port 4 e
rlabel m2 49 48 49 48 3 _clk
rlabel m2c 10 19 10 19 3 #7
rlabel m2c 10 45 10 45 3 CLK
port 4 e
rlabel m2 9 18 9 18 3 #7
rlabel m2 9 19 9 19 3 #7
rlabel m2 9 22 9 22 3 #7
rlabel m2 9 44 9 44 3 CLK
port 4 e
rlabel m2 9 45 9 45 3 CLK
port 4 e
rlabel m2 9 48 9 48 3 CLK
port 4 e
<< end >>
